
module huffman_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;

  ADDHXL U2 ( .A(A[6]), .B(n2), .CO(n1), .S(SUM[6]) );
  ADDHXL U3 ( .A(A[5]), .B(n3), .CO(n2), .S(SUM[5]) );
  ADDHXL U5 ( .A(A[3]), .B(n5), .CO(n4), .S(SUM[3]) );
  ADDHXL U6 ( .A(A[2]), .B(n6), .CO(n5), .S(SUM[2]) );
  ADDHXL U7 ( .A(A[1]), .B(A[0]), .CO(n6), .S(SUM[1]) );
  ADDHXL U4 ( .A(A[4]), .B(n4), .CO(n3), .S(SUM[4]) );
  INVX1 U11 ( .A(A[0]), .Y(SUM[0]) );
  AOI2BB2X1 U12 ( .B0(n1), .B1(A[7]), .A0N(n1), .A1N(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;

  ADDHXL U3 ( .A(A[5]), .B(n3), .CO(n2), .S(SUM[5]) );
  ADDHXL U4 ( .A(A[4]), .B(n4), .CO(n3), .S(SUM[4]) );
  ADDHXL U5 ( .A(A[3]), .B(n5), .CO(n4), .S(SUM[3]) );
  ADDHXL U2 ( .A(A[6]), .B(n2), .CO(n1), .S(SUM[6]) );
  ADDHXL U7 ( .A(A[1]), .B(A[0]), .CO(n6), .S(SUM[1]) );
  ADDHXL U6 ( .A(A[2]), .B(n6), .CO(n5), .S(SUM[2]) );
  AOI2BB2X1 U11 ( .B0(n1), .B1(A[7]), .A0N(n1), .A1N(A[7]), .Y(SUM[7]) );
  INVX1 U12 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module huffman_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;

  ADDHXL U2 ( .A(A[6]), .B(n2), .CO(n1), .S(SUM[6]) );
  ADDHXL U3 ( .A(A[5]), .B(n3), .CO(n2), .S(SUM[5]) );
  ADDHXL U4 ( .A(A[4]), .B(n4), .CO(n3), .S(SUM[4]) );
  ADDHXL U5 ( .A(A[3]), .B(n5), .CO(n4), .S(SUM[3]) );
  ADDHXL U6 ( .A(A[2]), .B(n6), .CO(n5), .S(SUM[2]) );
  ADDHXL U7 ( .A(A[1]), .B(A[0]), .CO(n6), .S(SUM[1]) );
  INVXL U11 ( .A(A[0]), .Y(SUM[0]) );
  AOI2BB2X1 U12 ( .B0(n1), .B1(A[7]), .A0N(n1), .A1N(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_3 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;

  ADDHXL U2 ( .A(A[6]), .B(n2), .CO(n1), .S(SUM[6]) );
  ADDHXL U3 ( .A(A[5]), .B(n3), .CO(n2), .S(SUM[5]) );
  ADDHXL U4 ( .A(A[4]), .B(n4), .CO(n3), .S(SUM[4]) );
  ADDHXL U5 ( .A(A[3]), .B(n5), .CO(n4), .S(SUM[3]) );
  ADDHXL U6 ( .A(A[2]), .B(n6), .CO(n5), .S(SUM[2]) );
  ADDHXL U7 ( .A(A[1]), .B(A[0]), .CO(n6), .S(SUM[1]) );
  INVX1 U11 ( .A(A[0]), .Y(SUM[0]) );
  AOI2BB2X1 U12 ( .B0(n1), .B1(A[7]), .A0N(n1), .A1N(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_4 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;

  ADDHXL U2 ( .A(A[6]), .B(n2), .CO(n1), .S(SUM[6]) );
  ADDHXL U3 ( .A(A[5]), .B(n3), .CO(n2), .S(SUM[5]) );
  ADDHXL U4 ( .A(A[4]), .B(n4), .CO(n3), .S(SUM[4]) );
  ADDHXL U5 ( .A(A[3]), .B(n5), .CO(n4), .S(SUM[3]) );
  ADDHXL U6 ( .A(A[2]), .B(n6), .CO(n5), .S(SUM[2]) );
  ADDHXL U7 ( .A(A[1]), .B(A[0]), .CO(n6), .S(SUM[1]) );
  AOI2BB2XL U11 ( .B0(n1), .B1(A[7]), .A0N(n1), .A1N(A[7]), .Y(SUM[7]) );
  INVX1 U12 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module huffman_DW01_inc_5 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;

  ADDHXL U2 ( .A(A[6]), .B(n2), .CO(n1), .S(SUM[6]) );
  ADDHXL U3 ( .A(A[5]), .B(n3), .CO(n2), .S(SUM[5]) );
  ADDHXL U4 ( .A(A[4]), .B(n4), .CO(n3), .S(SUM[4]) );
  ADDHXL U5 ( .A(A[3]), .B(n5), .CO(n4), .S(SUM[3]) );
  ADDHXL U6 ( .A(A[2]), .B(n6), .CO(n5), .S(SUM[2]) );
  ADDHXL U7 ( .A(A[1]), .B(A[0]), .CO(n6), .S(SUM[1]) );
  INVXL U11 ( .A(A[0]), .Y(SUM[0]) );
  AOI2BB2X1 U12 ( .B0(n1), .B1(A[7]), .A0N(n1), .A1N(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_add_2 ( A, B, CI, SUM, CO, IN0, IN1, IN2, IN3, IN4 );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI, IN0, IN1, IN2, IN3, IN4;
  output CO;
  wire   n5, n8, n11, n18, n20, n21, n22, n23, n24, n25, n26, n27, n28, n31,
         n32, n33, n34, n35, n36, n38, n39, n45, n46, n48, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n44, n107, n108, n109,
         n110, n111, n112, n113, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n139;
  assign n139 = IN0;

  NAND2X2 U15 ( .A(B[6]), .B(A[6]), .Y(n18) );
  NOR2X8 U30 ( .A(B[4]), .B(A[4]), .Y(n27) );
  NAND2X6 U63 ( .A(B[0]), .B(n80), .Y(n91) );
  CLKINVX6 U64 ( .A(n90), .Y(n80) );
  INVX1 U66 ( .A(n119), .Y(n48) );
  BUFX4 U68 ( .A(n39), .Y(n81) );
  NAND2X6 U70 ( .A(B[4]), .B(A[4]), .Y(n28) );
  NOR2X8 U74 ( .A(B[2]), .B(A[2]), .Y(n34) );
  NAND2X6 U76 ( .A(B[2]), .B(A[2]), .Y(n35) );
  CLKINVX1 U77 ( .A(A[0]), .Y(n90) );
  CLKINVX3 U81 ( .A(n31), .Y(n46) );
  AND2X2 U83 ( .A(n133), .B(n89), .Y(SUM[0]) );
  INVX3 U84 ( .A(n34), .Y(n93) );
  OR2XL U91 ( .A(B[0]), .B(A[0]), .Y(n103) );
  OAI21X4 U94 ( .A0(n38), .A1(n91), .B0(n39), .Y(n102) );
  OR2X8 U103 ( .A(B[6]), .B(A[6]), .Y(n104) );
  NOR2X8 U106 ( .A(B[3]), .B(A[3]), .Y(n31) );
  NAND2X4 U108 ( .A(A[3]), .B(B[3]), .Y(n32) );
  NAND2X4 U109 ( .A(A[1]), .B(B[1]), .Y(n39) );
  INVX1 U113 ( .A(n22), .Y(n20) );
  CLKINVX1 U115 ( .A(n27), .Y(n45) );
  DFFSX1 R_298 ( .D(n103), .CK(n139), .SN(IN1), .Q(n133) );
  DFFSX1 R_305 ( .D(n38), .CK(n139), .SN(IN1), .Q(n132) );
  DFFSX1 R_307 ( .D(n39), .CK(n139), .SN(IN1), .Q(n131) );
  DFFRX1 R_315 ( .D(n101), .CK(n139), .RN(IN2), .Q(n129) );
  DFFSX1 R_314 ( .D(n102), .CK(n139), .SN(IN2), .Q(n130) );
  DFFSX1 R_319 ( .D(n46), .CK(n139), .SN(IN1), .Q(n128) );
  DFFRX1 R_320 ( .D(n32), .CK(n139), .RN(IN1), .Q(n127) );
  DFFSX1 R_345 ( .D(n18), .CK(n139), .SN(IN1), .Q(n126) );
  NAND2X1 U5 ( .A(IN4), .B(n123), .Y(n11) );
  NAND2X4 U73 ( .A(B[5]), .B(A[5]), .Y(n25) );
  NOR2X8 U71 ( .A(B[5]), .B(A[5]), .Y(n24) );
  NOR2X6 U110 ( .A(B[1]), .B(A[1]), .Y(n38) );
  DFFRX1 R_200_RW ( .D(n35), .CK(n139), .RN(IN1), .Q(n135) );
  NOR2X6 U111 ( .A(n31), .B(n34), .Y(n101) );
  DFFSX1 R_368 ( .D(n81), .CK(n139), .SN(IN1), .Q(n125) );
  DFFSX1 R_370 ( .D(n45), .CK(n139), .SN(IN1), .Q(n124) );
  DFFSX1 R_389 ( .D(n31), .CK(n139), .SN(IN2), .Q(n122) );
  DFFSX1 R_390 ( .D(n32), .CK(n139), .SN(IN2), .Q(n121) );
  DFFSX1 R_288 ( .D(n25), .CK(n139), .SN(IN3), .Q(n134) );
  DFFRX1 R_396 ( .D(n24), .CK(n139), .RN(IN3), .Q(n120) );
  DFFSX1 R_407 ( .D(A[7]), .CK(n139), .SN(IN2), .Q(n118) );
  DFFSX1 R_427 ( .D(n28), .CK(n139), .SN(IN1), .Q(n117) );
  DFFRX1 R_428 ( .D(n25), .CK(n139), .RN(IN1), .Q(n116) );
  DFFRX1 R_429 ( .D(n18), .CK(n139), .RN(IN2), .Q(n115) );
  DFFRX1 R_400_RW ( .D(n38), .CK(n139), .RN(IN1), .Q(n119) );
  DFFSX1 R_444 ( .D(n104), .CK(n139), .SN(IN2), .Q(n113) );
  DFFSX1 R_453 ( .D(n27), .CK(n139), .SN(IN2), .Q(n112) );
  DFFSX1 R_454 ( .D(n91), .CK(n139), .SN(IN1), .Q(n111) );
  DFFRX1 R_455 ( .D(n28), .CK(n139), .RN(IN1), .Q(n110) );
  DFFSX1 R_456 ( .D(n35), .CK(n139), .SN(IN2), .Q(n109) );
  DFFSX1 R_457 ( .D(n93), .CK(n139), .SN(IN1), .Q(n108) );
  DFFSX1 R_458 ( .D(n24), .CK(n139), .SN(IN1), .Q(n107) );
  DFFRXL R_387 ( .D(A[7]), .CK(n139), .RN(IN2), .Q(n123) );
  CLKBUFX3 U61 ( .A(n111), .Y(n89) );
  CLKINVX1 U62 ( .A(n115), .Y(n98) );
  OAI21XL U65 ( .A0(n107), .A1(n117), .B0(n116), .Y(n23) );
  NOR2X1 U67 ( .A(n107), .B(n112), .Y(n22) );
  OR2X1 U69 ( .A(IN4), .B(n118), .Y(n105) );
  NAND2X1 U72 ( .A(n22), .B(n113), .Y(n99) );
  CLKBUFX3 U75 ( .A(n120), .Y(n82) );
  CLKINVX1 U78 ( .A(n82), .Y(n44) );
  AND2X2 U79 ( .A(n44), .B(n134), .Y(n84) );
  OAI21XL U80 ( .A0(n109), .A1(n122), .B0(n121), .Y(n100) );
  NAND2X1 U82 ( .A(n108), .B(n109), .Y(n92) );
  NAND2X1 U85 ( .A(n124), .B(n110), .Y(n5) );
  NAND2X1 U86 ( .A(n125), .B(n48), .Y(n8) );
  AND2X2 U87 ( .A(n113), .B(n126), .Y(n85) );
  AND2X2 U88 ( .A(n128), .B(n127), .Y(n87) );
  AND2X2 U89 ( .A(n130), .B(n129), .Y(n94) );
  OAI21XL U90 ( .A0(n132), .A1(n111), .B0(n131), .Y(n83) );
  CLKINVX1 U92 ( .A(n23), .Y(n21) );
  CLKINVX1 U93 ( .A(n83), .Y(n36) );
  NOR2X1 U95 ( .A(n94), .B(n100), .Y(n95) );
  AOI21X1 U96 ( .A0(n113), .A1(n23), .B0(n98), .Y(n97) );
  AND2X2 U97 ( .A(n105), .B(n11), .Y(n86) );
  XOR2X1 U98 ( .A(n8), .B(n89), .Y(SUM[1]) );
  OAI2BB1X1 U99 ( .A0N(n108), .A1N(n83), .B0(n135), .Y(n33) );
  OAI21XL U100 ( .A0(n95), .A1(n99), .B0(n97), .Y(n96) );
  OAI21XL U101 ( .A0(n95), .A1(n20), .B0(n21), .Y(n88) );
  OAI21XL U102 ( .A0(n95), .A1(n112), .B0(n110), .Y(n26) );
  XOR2X1 U104 ( .A(n36), .B(n92), .Y(SUM[2]) );
  XOR2X1 U105 ( .A(n33), .B(n87), .Y(SUM[3]) );
  XOR2X1 U107 ( .A(n26), .B(n84), .Y(SUM[5]) );
  XOR2X1 U112 ( .A(n95), .B(n5), .Y(SUM[4]) );
  XOR2X1 U114 ( .A(n96), .B(n86), .Y(SUM[7]) );
  XOR2X1 U116 ( .A(n88), .B(n85), .Y(SUM[6]) );
endmodule


module huffman_add_314_DP_OP_292_9816_0 ( I1, I2, O2 );
  input [7:0] I1;
  input [7:0] I2;
  output [7:0] O2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36;
  assign O2[0] = n13;
  assign O2[1] = n14;
  assign O2[2] = n15;
  assign O2[3] = n16;
  assign O2[4] = n17;
  assign O2[5] = n18;
  assign O2[6] = n19;
  assign O2[7] = n20;
  assign n21 = I2[0];
  assign n22 = I2[1];
  assign n23 = I2[2];
  assign n24 = I2[3];
  assign n25 = I2[4];
  assign n26 = I2[5];
  assign n27 = I2[6];
  assign n28 = I2[7];
  assign n29 = I1[0];
  assign n30 = I1[1];
  assign n31 = I1[2];
  assign n32 = I1[3];
  assign n33 = I1[4];
  assign n34 = I1[5];
  assign n35 = I1[6];
  assign n36 = I1[7];

  ADDFXL U3 ( .A(n35), .B(n27), .CI(n3), .CO(n2), .S(n19) );
  ADDFXL U4 ( .A(n34), .B(n26), .CI(n4), .CO(n3), .S(n18) );
  ADDFXL U5 ( .A(n33), .B(n25), .CI(n5), .CO(n4), .S(n17) );
  ADDFXL U6 ( .A(n32), .B(n24), .CI(n6), .CO(n5), .S(n16) );
  ADDFXL U7 ( .A(n31), .B(n23), .CI(n7), .CO(n6), .S(n15) );
  ADDFXL U8 ( .A(n30), .B(n22), .CI(n8), .CO(n7), .S(n14) );
  ADDHXL U9 ( .A(n21), .B(n29), .CO(n8), .S(n13) );
  XOR2X1 U2 ( .A(n36), .B(n28), .Y(n1) );
  XOR2X1 U1 ( .A(n2), .B(n1), .Y(n20) );
endmodule


module huffman_add_318_DP_OP_291_9816_1 ( I1, I2, O1, IN0, IN1, IN2 );
  input [7:0] I1;
  input [7:0] I2;
  output [7:0] O1;
  input IN0, IN1, IN2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n11, n12, n14, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n41, n44, n45, n46, n47, n48, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n88,
         n89, n90, n91, n92, n93, n95, n96, n98, n99;
  assign O1[1] = n55;
  assign O1[2] = n56;
  assign O1[3] = n57;
  assign O1[4] = n58;
  assign O1[5] = n59;
  assign O1[6] = n60;
  assign O1[7] = n61;
  assign n62 = I2[0];
  assign n63 = I2[1];
  assign n64 = I2[2];
  assign n65 = I2[3];
  assign n66 = I2[4];
  assign n67 = I2[5];
  assign n68 = I2[6];
  assign n69 = I2[7];
  assign n70 = I1[0];
  assign n71 = I1[1];
  assign n72 = I1[2];
  assign n73 = I1[3];
  assign n74 = I1[4];
  assign n75 = I1[5];
  assign n76 = I1[6];
  assign n77 = I1[7];
  assign n98 = IN0;

  AOI21X1 U9 ( .A0(n23), .A1(n83), .B0(n16), .Y(n14) );
  NAND2X1 U5 ( .A(n69), .B(n77), .Y(n11) );
  NAND2X2 U52 ( .A(n63), .B(n71), .Y(n39) );
  NOR2X2 U38 ( .A(n65), .B(n73), .Y(n31) );
  NAND2X2 U31 ( .A(n66), .B(n74), .Y(n28) );
  NAND2X1 U15 ( .A(n68), .B(n76), .Y(n18) );
  NAND2X1 U2 ( .A(n84), .B(n11), .Y(n2) );
  NAND2X1 U28 ( .A(n45), .B(n28), .Y(n5) );
  XOR2X1 U26 ( .A(n88), .B(n87), .Y(n58) );
  NAND2X1 U42 ( .A(n47), .B(n35), .Y(n7) );
  XOR2X1 U40 ( .A(n36), .B(n7), .Y(n56) );
  NAND2X1 U22 ( .A(n44), .B(n25), .Y(n4) );
  NAND2X1 U36 ( .A(n46), .B(n32), .Y(n6) );
  NAND2X1 U12 ( .A(n83), .B(n18), .Y(n3) );
  NAND2X1 U49 ( .A(n48), .B(n39), .Y(n8) );
  XOR2X1 U46 ( .A(n8), .B(n41), .Y(n55) );
  OAI21X4 U21 ( .A0(n24), .A1(n28), .B0(n25), .Y(n23) );
  INVX2 U61 ( .A(n1), .Y(n79) );
  NOR2X4 U62 ( .A(n24), .B(n27), .Y(n22) );
  CLKAND2X3 U63 ( .A(n22), .B(n83), .Y(n78) );
  OAI21X2 U65 ( .A0(n36), .A1(n34), .B0(n35), .Y(n33) );
  OAI21X4 U66 ( .A0(n1), .A1(n27), .B0(n28), .Y(n26) );
  NOR2X8 U67 ( .A(n67), .B(n75), .Y(n24) );
  OAI2BB1X4 U68 ( .A0N(n78), .A1N(n79), .B0(n14), .Y(n12) );
  AND2X8 U69 ( .A(n82), .B(n80), .Y(n1) );
  NAND2X4 U70 ( .A(n81), .B(n37), .Y(n80) );
  OAI21X4 U71 ( .A0(n38), .A1(n41), .B0(n39), .Y(n37) );
  NAND2X4 U72 ( .A(n62), .B(n70), .Y(n41) );
  NOR2X6 U73 ( .A(n63), .B(n71), .Y(n38) );
  NOR2X6 U75 ( .A(n64), .B(n72), .Y(n34) );
  OA21X4 U76 ( .A0(n31), .A1(n35), .B0(n32), .Y(n82) );
  NAND2X4 U77 ( .A(n64), .B(n72), .Y(n35) );
  OAI21X4 U79 ( .A0(n1), .A1(n20), .B0(n21), .Y(n19) );
  NAND2X4 U80 ( .A(n67), .B(n75), .Y(n25) );
  NOR2X4 U81 ( .A(n66), .B(n74), .Y(n27) );
  CLKINVX1 U82 ( .A(n38), .Y(n48) );
  INVX1 U83 ( .A(n23), .Y(n21) );
  INVX1 U84 ( .A(n22), .Y(n20) );
  INVX1 U85 ( .A(n31), .Y(n46) );
  INVX1 U86 ( .A(n24), .Y(n44) );
  CLKINVX1 U87 ( .A(n34), .Y(n47) );
  INVX3 U88 ( .A(n37), .Y(n36) );
  INVX1 U89 ( .A(n27), .Y(n45) );
  OR2X1 U90 ( .A(n69), .B(n77), .Y(n84) );
  INVX1 U91 ( .A(n18), .Y(n16) );
  CLKAND2X3 U93 ( .A(n85), .B(n41), .Y(O1[0]) );
  OR2X2 U94 ( .A(n62), .B(n70), .Y(n85) );
  DFFSX1 R_321 ( .D(n12), .CK(n98), .SN(IN1), .Q(n99) );
  DFFSX1 R_322 ( .D(n2), .CK(n98), .SN(IN1), .Q(n96) );
  OR2X2 U92 ( .A(n68), .B(n76), .Y(n83) );
  NAND2X4 U60 ( .A(n65), .B(n73), .Y(n32) );
  NOR2X6 U74 ( .A(n31), .B(n34), .Y(n81) );
  DFFSX1 R_364 ( .D(n26), .CK(n98), .SN(IN2), .Q(n95) );
  DFFRX1 R_365 ( .D(n4), .CK(n98), .RN(IN2), .Q(n93) );
  DFFSX1 R_366 ( .D(n19), .CK(n98), .SN(IN2), .Q(n92) );
  DFFRX1 R_367 ( .D(n3), .CK(n98), .RN(IN2), .Q(n91) );
  DFFSX1 R_374 ( .D(n33), .CK(n98), .SN(IN2), .Q(n90) );
  DFFRX1 R_375 ( .D(n6), .CK(n98), .RN(IN2), .Q(n89) );
  DFFSX1 R_377 ( .D(n1), .CK(n98), .SN(IN2), .Q(n88) );
  DFFSX1 R_378 ( .D(n5), .CK(n98), .SN(IN2), .Q(n87) );
  XNOR2X1 U64 ( .A(n90), .B(n89), .Y(n57) );
  XNOR2X1 U78 ( .A(n92), .B(n91), .Y(n60) );
  XNOR2X1 U95 ( .A(n95), .B(n93), .Y(n59) );
  XNOR2X1 U96 ( .A(n99), .B(n96), .Y(n61) );
endmodule


module huffman_add_303_DP_OP_294_9816_1 ( I1, I2, O2, IN0, IN1, IN2, IN3 );
  input [7:0] I1;
  input [7:0] I2;
  output [7:0] O2;
  input IN0, IN1, IN2, IN3;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n11, n12, n13, n14, n16, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n41, n45, n46, n47, n48, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n92, n94, n95, n96, n98;
  assign O2[1] = n55;
  assign O2[2] = n56;
  assign O2[3] = n57;
  assign O2[4] = n58;
  assign O2[5] = n59;
  assign O2[6] = n60;
  assign O2[7] = n61;
  assign n62 = I2[0];
  assign n63 = I2[1];
  assign n64 = I2[2];
  assign n65 = I2[3];
  assign n66 = I2[4];
  assign n67 = I2[5];
  assign n68 = I2[6];
  assign n69 = I2[7];
  assign n70 = I1[0];
  assign n71 = I1[1];
  assign n72 = I1[2];
  assign n73 = I1[3];
  assign n74 = I1[4];
  assign n75 = I1[5];
  assign n76 = I1[6];
  assign n77 = I1[7];
  assign n98 = IN0;

  NAND2X1 U5 ( .A(n77), .B(n69), .Y(n11) );
  AOI21X4 U33 ( .A0(n37), .A1(n29), .B0(n30), .Y(n1) );
  NAND2X2 U57 ( .A(n70), .B(n62), .Y(n41) );
  NAND2X1 U52 ( .A(n71), .B(n63), .Y(n39) );
  NOR2X2 U44 ( .A(n72), .B(n64), .Y(n34) );
  NAND2X1 U42 ( .A(n47), .B(n35), .Y(n7) );
  XOR2X1 U40 ( .A(n36), .B(n7), .Y(n56) );
  NOR2X1 U34 ( .A(n34), .B(n31), .Y(n29) );
  NAND2X1 U39 ( .A(n73), .B(n65), .Y(n32) );
  OAI21X1 U35 ( .A0(n31), .A1(n35), .B0(n32), .Y(n30) );
  NOR2X2 U30 ( .A(n74), .B(n66), .Y(n27) );
  NAND2X2 U31 ( .A(n74), .B(n66), .Y(n28) );
  NAND2X1 U28 ( .A(n45), .B(n28), .Y(n5) );
  XOR2X1 U26 ( .A(n83), .B(n90), .Y(n58) );
  NAND2X1 U49 ( .A(n48), .B(n39), .Y(n8) );
  XOR2X1 U46 ( .A(n8), .B(n41), .Y(n55) );
  NAND2X1 U36 ( .A(n46), .B(n32), .Y(n6) );
  XNOR2X1 U32 ( .A(n89), .B(n88), .Y(n57) );
  NOR2X2 U24 ( .A(n75), .B(n67), .Y(n24) );
  NAND2X1 U22 ( .A(n78), .B(n25), .Y(n4) );
  NAND2X1 U15 ( .A(n76), .B(n68), .Y(n18) );
  AOI21X1 U9 ( .A0(n23), .A1(n80), .B0(n16), .Y(n14) );
  NAND2X1 U2 ( .A(n81), .B(n11), .Y(n2) );
  NAND2X1 U12 ( .A(n80), .B(n18), .Y(n3) );
  OAI21X4 U41 ( .A0(n36), .A1(n34), .B0(n35), .Y(n33) );
  NOR2X4 U60 ( .A(n73), .B(n65), .Y(n31) );
  INVX3 U61 ( .A(n23), .Y(n21) );
  NAND2X6 U62 ( .A(n72), .B(n64), .Y(n35) );
  OAI21X2 U63 ( .A0(n1), .A1(n13), .B0(n14), .Y(n12) );
  OAI21X4 U64 ( .A0(n24), .A1(n28), .B0(n25), .Y(n23) );
  NAND2X2 U65 ( .A(n22), .B(n80), .Y(n13) );
  NOR2X2 U66 ( .A(n27), .B(n24), .Y(n22) );
  NAND2X4 U68 ( .A(n75), .B(n67), .Y(n25) );
  OAI21X4 U69 ( .A0(n38), .A1(n41), .B0(n39), .Y(n37) );
  NOR2X4 U70 ( .A(n71), .B(n63), .Y(n38) );
  OR2X4 U71 ( .A(n75), .B(n67), .Y(n78) );
  INVX1 U72 ( .A(n22), .Y(n20) );
  OR2X1 U73 ( .A(n77), .B(n69), .Y(n81) );
  INVX1 U74 ( .A(n18), .Y(n16) );
  OR2X2 U75 ( .A(n76), .B(n68), .Y(n80) );
  INVX1 U76 ( .A(n31), .Y(n46) );
  CLKAND2X3 U77 ( .A(n82), .B(n41), .Y(O2[0]) );
  OR2X1 U78 ( .A(n70), .B(n62), .Y(n82) );
  INVX1 U79 ( .A(n38), .Y(n48) );
  INVX1 U80 ( .A(n27), .Y(n45) );
  INVX1 U81 ( .A(n34), .Y(n47) );
  INVX3 U82 ( .A(n37), .Y(n36) );
  DFFSX1 R_197_RW ( .D(n3), .CK(n98), .SN(IN1), .Q(n96) );
  DFFSX1 R_260 ( .D(n4), .CK(n98), .SN(IN1), .Q(n95) );
  DFFSX1 R_261 ( .D(n12), .CK(n98), .SN(IN2), .Q(n94) );
  DFFSX1 R_262 ( .D(n2), .CK(n98), .SN(IN2), .Q(n92) );
  DFFRX1 R_313 ( .D(n5), .CK(n98), .RN(IN3), .Q(n90) );
  DFFSX1 R_327 ( .D(n33), .CK(n98), .SN(IN3), .Q(n89) );
  DFFSX1 R_328_RW ( .D(n6), .CK(n98), .SN(IN2), .Q(n88) );
  DFFSX1 R_419 ( .D(n27), .CK(n98), .SN(IN1), .Q(n87) );
  DFFRX1 R_420 ( .D(n28), .CK(n98), .RN(IN1), .Q(n86) );
  DFFSX1 R_434 ( .D(n20), .CK(n98), .SN(IN1), .Q(n85) );
  DFFRX1 R_435 ( .D(n21), .CK(n98), .RN(IN1), .Q(n84) );
  DFFSX1 R_445 ( .D(n1), .CK(n98), .SN(IN1), .Q(n83) );
  OAI21XL U67 ( .A0(n83), .A1(n85), .B0(n84), .Y(n19) );
  OAI21XL U83 ( .A0(n83), .A1(n87), .B0(n86), .Y(n26) );
  XNOR2X1 U84 ( .A(n94), .B(n92), .Y(n61) );
  XNOR2X1 U85 ( .A(n26), .B(n95), .Y(n59) );
  XNOR2X1 U86 ( .A(n19), .B(n96), .Y(n60) );
endmodule


module huffman_add_307_DP_OP_293_9816_1 ( I1, I2, O1 );
  input [7:0] I1;
  input [7:0] I2;
  output [7:0] O1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n11, n12, n13, n14, n16, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n41, n44, n45, n46, n47, n48, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80;
  assign O1[1] = n55;
  assign O1[2] = n56;
  assign O1[3] = n57;
  assign O1[4] = n58;
  assign O1[5] = n59;
  assign O1[6] = n60;
  assign O1[7] = n61;
  assign n62 = I2[0];
  assign n63 = I2[1];
  assign n64 = I2[2];
  assign n65 = I2[3];
  assign n66 = I2[4];
  assign n67 = I2[5];
  assign n68 = I2[6];
  assign n69 = I2[7];
  assign n70 = I1[0];
  assign n71 = I1[1];
  assign n72 = I1[2];
  assign n73 = I1[3];
  assign n74 = I1[4];
  assign n75 = I1[5];
  assign n76 = I1[6];
  assign n77 = I1[7];

  NAND2X1 U8 ( .A(n22), .B(n78), .Y(n13) );
  NAND2X1 U15 ( .A(n68), .B(n76), .Y(n18) );
  AOI21X1 U9 ( .A0(n23), .A1(n78), .B0(n16), .Y(n14) );
  NAND2X1 U5 ( .A(n69), .B(n77), .Y(n11) );
  NAND2X1 U2 ( .A(n79), .B(n11), .Y(n2) );
  NAND2X2 U45 ( .A(n64), .B(n72), .Y(n35) );
  OAI21X1 U21 ( .A0(n24), .A1(n28), .B0(n25), .Y(n23) );
  NOR2X1 U51 ( .A(n63), .B(n71), .Y(n38) );
  NAND2X2 U57 ( .A(n62), .B(n70), .Y(n41) );
  NAND2X1 U52 ( .A(n63), .B(n71), .Y(n39) );
  NOR2X2 U44 ( .A(n64), .B(n72), .Y(n34) );
  NAND2X1 U42 ( .A(n47), .B(n35), .Y(n7) );
  XOR2X1 U40 ( .A(n36), .B(n7), .Y(n56) );
  NOR2X2 U38 ( .A(n65), .B(n73), .Y(n31) );
  NOR2X1 U34 ( .A(n31), .B(n34), .Y(n29) );
  NAND2X1 U39 ( .A(n65), .B(n73), .Y(n32) );
  OAI21X1 U35 ( .A0(n31), .A1(n35), .B0(n32), .Y(n30) );
  NOR2X2 U30 ( .A(n66), .B(n74), .Y(n27) );
  NAND2X2 U31 ( .A(n66), .B(n74), .Y(n28) );
  NAND2X1 U28 ( .A(n45), .B(n28), .Y(n5) );
  XOR2X1 U26 ( .A(n1), .B(n5), .Y(n58) );
  NAND2X1 U49 ( .A(n48), .B(n39), .Y(n8) );
  XOR2X1 U46 ( .A(n8), .B(n41), .Y(n55) );
  OAI21X1 U41 ( .A0(n36), .A1(n34), .B0(n35), .Y(n33) );
  NAND2X1 U36 ( .A(n46), .B(n32), .Y(n6) );
  XNOR2X1 U32 ( .A(n33), .B(n6), .Y(n57) );
  OAI21X1 U27 ( .A0(n1), .A1(n27), .B0(n28), .Y(n26) );
  NOR2X2 U24 ( .A(n67), .B(n75), .Y(n24) );
  NAND2X1 U25 ( .A(n67), .B(n75), .Y(n25) );
  NAND2X1 U22 ( .A(n44), .B(n25), .Y(n4) );
  XNOR2X1 U16 ( .A(n26), .B(n4), .Y(n59) );
  NOR2X1 U20 ( .A(n27), .B(n24), .Y(n22) );
  XNOR2X1 U1 ( .A(n12), .B(n2), .Y(n61) );
  NAND2X1 U12 ( .A(n78), .B(n18), .Y(n3) );
  XNOR2X1 U6 ( .A(n19), .B(n3), .Y(n60) );
  OAI21X2 U60 ( .A0(n1), .A1(n20), .B0(n21), .Y(n19) );
  AOI21X4 U61 ( .A0(n37), .A1(n29), .B0(n30), .Y(n1) );
  INVX2 U62 ( .A(n37), .Y(n36) );
  OAI21X4 U63 ( .A0(n38), .A1(n41), .B0(n39), .Y(n37) );
  OAI21X2 U64 ( .A0(n1), .A1(n13), .B0(n14), .Y(n12) );
  INVX1 U65 ( .A(n18), .Y(n16) );
  OR2X1 U66 ( .A(n68), .B(n76), .Y(n78) );
  INVX1 U67 ( .A(n24), .Y(n44) );
  INVX1 U68 ( .A(n31), .Y(n46) );
  AND2X2 U69 ( .A(n80), .B(n41), .Y(O1[0]) );
  OR2X1 U70 ( .A(n62), .B(n70), .Y(n80) );
  INVX1 U71 ( .A(n38), .Y(n48) );
  INVX1 U72 ( .A(n27), .Y(n45) );
  INVX1 U73 ( .A(n34), .Y(n47) );
  INVX1 U74 ( .A(n23), .Y(n21) );
  INVX1 U75 ( .A(n22), .Y(n20) );
  OR2X1 U76 ( .A(n69), .B(n77), .Y(n79) );
endmodule


module huffman_DW01_add_13 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n10, n11, n12, n13, n14, n16, n18, n19,
         n20, n21, n22, n24, n26, n27, n28, n29, n30, n32, n34, n35, n37, n39,
         n41, n43, n76, n77, n78, n79, n80, n81;

  NAND2X1 U11 ( .A(B[6]), .B(A[6]), .Y(n13) );
  NAND2X1 U5 ( .A(B[7]), .B(A[7]), .Y(n10) );
  NAND2X1 U2 ( .A(n81), .B(n10), .Y(n1) );
  XNOR2X1 U1 ( .A(n11), .B(n1), .Y(SUM[7]) );
  NAND2X1 U8 ( .A(n39), .B(n13), .Y(n2) );
  XOR2X1 U6 ( .A(n14), .B(n2), .Y(SUM[6]) );
  NAND2X1 U16 ( .A(n79), .B(n18), .Y(n3) );
  XNOR2X1 U12 ( .A(n19), .B(n3), .Y(SUM[5]) );
  NAND2X1 U22 ( .A(n41), .B(n21), .Y(n4) );
  XOR2X1 U20 ( .A(n22), .B(n4), .Y(SUM[4]) );
  NAND2X1 U30 ( .A(n77), .B(n26), .Y(n5) );
  XNOR2X1 U26 ( .A(n27), .B(n5), .Y(SUM[3]) );
  NAND2X1 U36 ( .A(n43), .B(n29), .Y(n6) );
  XOR2X1 U34 ( .A(n30), .B(n6), .Y(SUM[2]) );
  XNOR2X1 U40 ( .A(n7), .B(n35), .Y(SUM[1]) );
  OAI21X1 U7 ( .A0(n14), .A1(n12), .B0(n13), .Y(n11) );
  AOI21X2 U41 ( .A0(n78), .A1(n35), .B0(n32), .Y(n30) );
  OAI21X2 U35 ( .A0(n30), .A1(n28), .B0(n29), .Y(n27) );
  AOI21X2 U27 ( .A0(n27), .A1(n77), .B0(n24), .Y(n22) );
  OAI21X2 U21 ( .A0(n22), .A1(n20), .B0(n21), .Y(n19) );
  AOI21X2 U13 ( .A0(n19), .A1(n79), .B0(n16), .Y(n14) );
  NAND2X1 U19 ( .A(B[5]), .B(A[5]), .Y(n18) );
  NAND2X1 U44 ( .A(n78), .B(n34), .Y(n7) );
  CLKINVX1 U57 ( .A(n37), .Y(n35) );
  NAND2X1 U58 ( .A(B[0]), .B(A[0]), .Y(n37) );
  NOR2X1 U59 ( .A(n76), .B(A[4]), .Y(n20) );
  NOR2X1 U60 ( .A(B[6]), .B(A[6]), .Y(n12) );
  OR2XL U61 ( .A(B[5]), .B(A[5]), .Y(n79) );
  NAND2X1 U62 ( .A(n76), .B(A[4]), .Y(n21) );
  NAND2X1 U63 ( .A(B[3]), .B(A[3]), .Y(n26) );
  OR2X1 U64 ( .A(B[3]), .B(A[3]), .Y(n77) );
  AND2X2 U65 ( .A(n80), .B(n37), .Y(SUM[0]) );
  OR2XL U66 ( .A(B[0]), .B(A[0]), .Y(n80) );
  CLKBUFX2 U67 ( .A(B[4]), .Y(n76) );
  NOR2XL U68 ( .A(B[2]), .B(A[2]), .Y(n28) );
  NAND2XL U69 ( .A(B[2]), .B(A[2]), .Y(n29) );
  NAND2X1 U70 ( .A(B[1]), .B(A[1]), .Y(n34) );
  OR2X1 U71 ( .A(B[1]), .B(A[1]), .Y(n78) );
  INVX1 U72 ( .A(n28), .Y(n43) );
  INVX1 U73 ( .A(n12), .Y(n39) );
  CLKINVX1 U74 ( .A(n20), .Y(n41) );
  CLKINVX1 U75 ( .A(n18), .Y(n16) );
  CLKINVX1 U76 ( .A(n26), .Y(n24) );
  CLKINVX1 U77 ( .A(n34), .Y(n32) );
  OR2X1 U78 ( .A(B[7]), .B(A[7]), .Y(n81) );
endmodule


module huffman ( clk, reset, gray_data, gray_valid, CNT_valid, CNT1, CNT2, 
        CNT3, CNT4, CNT5, CNT6, code_valid, HC1, HC2, HC3, HC4, HC5, HC6, M1, 
        M2, M3, M4, M5, M6 );
  input [7:0] gray_data;
  output [7:0] CNT1;
  output [7:0] CNT2;
  output [7:0] CNT3;
  output [7:0] CNT4;
  output [7:0] CNT5;
  output [7:0] CNT6;
  output [7:0] HC1;
  output [7:0] HC2;
  output [7:0] HC3;
  output [7:0] HC4;
  output [7:0] HC5;
  output [7:0] HC6;
  output [7:0] M1;
  output [7:0] M2;
  output [7:0] M3;
  output [7:0] M4;
  output [7:0] M5;
  output [7:0] M6;
  input clk, reset, gray_valid;
  output CNT_valid, code_valid;
  wire   re_order_en, out_en, N202, N203, N204, N205, N644, N645, N646, N647,
         N648, N649, N650, N651, N652, N653, N654, N658, N659, N660, N661,
         N662, N663, N664, N665, N666, N667, N668, N672, N673, N674, N675,
         N676, N677, N678, N679, N680, N681, N682, N686, N687, N688, N689,
         N690, N691, N692, N693, N694, N695, N696, N700, N701, N702, N703,
         N704, N705, N706, N707, N708, N709, N710, N714, N715, N716, N717,
         N718, N719, N720, N721, N722, N723, N724, N766, N767, N768, N769,
         N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780,
         N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791,
         N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802,
         N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813,
         \com[0][7] , \com[0][6] , \com[0][5] , \com[0][4] , \com[0][3] ,
         \com[0][2] , \com[0][1] , \com[0][0] , \com[1][7] , \com[1][6] ,
         \com[1][5] , \com[1][4] , \com[1][3] , \com[1][2] , \com[1][1] ,
         \com[1][0] , \com[2][7] , \com[2][6] , \com[2][5] , \com[2][4] ,
         \com[2][3] , \com[2][2] , \com[2][1] , \com[2][0] , \com[3][7] ,
         \com[3][6] , \com[3][5] , \com[3][4] , \com[3][3] , \com[3][1] ,
         \com[3][0] , \com[4][7] , \com[4][6] , \com[4][5] , \com[4][4] ,
         \com[4][3] , \com[4][2] , \com[4][1] , \com[4][0] , N1140, N1141,
         N1142, N1143, N1144, N1145, N1146, N1147, N1215, N1216, N1217, N1218,
         N1219, N1220, N1221, N1222, n474, n475, n477, n479, n481, n483, n485,
         n491, n493, n495, n497, n505, n507, n509, n511, n520, n522, n524,
         n526, n529, n531, n533, n535, n538, n540, n542, n544, n547, n549,
         n551, n553, n579, n605, n606, n607, n608, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n647, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n690, n691, n692, n693, n694, n695, n696, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n716, n717, n718, n719, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1198, n1199, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1766, n1767, n1768, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n2455, n2469,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254;
  wire   [2:0] state;
  wire   [2:0] next_state;
  wire   [7:0] com_after_1;
  wire   [2:0] tree_mem;
  wire   [2:0] tree_mem_back;
  assign HC1[7] = 1'b0;
  assign HC1[6] = 1'b0;
  assign HC1[5] = 1'b0;
  assign HC2[7] = 1'b0;
  assign HC2[6] = 1'b0;
  assign HC2[5] = 1'b0;
  assign HC3[7] = 1'b0;
  assign HC3[6] = 1'b0;
  assign HC3[5] = 1'b0;
  assign HC4[7] = 1'b0;
  assign HC4[6] = 1'b0;
  assign HC4[5] = 1'b0;
  assign HC5[7] = 1'b0;
  assign HC5[6] = 1'b0;
  assign HC5[5] = 1'b0;
  assign HC6[7] = 1'b0;
  assign HC6[6] = 1'b0;
  assign HC6[5] = 1'b0;
  assign M1[7] = 1'b0;
  assign M1[6] = 1'b0;
  assign M1[5] = 1'b0;
  assign M2[7] = 1'b0;
  assign M2[6] = 1'b0;
  assign M2[5] = 1'b0;
  assign M3[7] = 1'b0;
  assign M3[6] = 1'b0;
  assign M3[5] = 1'b0;
  assign M4[7] = 1'b0;
  assign M4[6] = 1'b0;
  assign M4[5] = 1'b0;
  assign M5[7] = 1'b0;
  assign M5[6] = 1'b0;
  assign M5[5] = 1'b0;
  assign M6[7] = 1'b0;
  assign M6[6] = 1'b0;
  assign M6[5] = 1'b0;

  DFFRX4 \CNT4_reg[2]  ( .D(n863), .CK(clk), .RN(n1804), .Q(CNT4[2]), .QN(n677) );
  DFFRX4 \CNT4_reg[3]  ( .D(n862), .CK(clk), .RN(n1804), .Q(CNT4[3]), .QN(n676) );
  DFFRX4 \CNT4_reg[4]  ( .D(n861), .CK(clk), .RN(n1811), .Q(CNT4[4]), .QN(n675) );
  DFFRX4 \CNT4_reg[7]  ( .D(n858), .CK(clk), .RN(n1811), .Q(CNT4[7]), .QN(n672) );
  DFFRX4 \CNT3_reg[1]  ( .D(n848), .CK(clk), .RN(n1813), .Q(CNT3[1]), .QN(n662) );
  DFFRX4 \CNT3_reg[2]  ( .D(n847), .CK(clk), .RN(n1813), .Q(CNT3[2]), .QN(n661) );
  DFFRX4 \CNT3_reg[3]  ( .D(n846), .CK(clk), .RN(n1813), .Q(CNT3[3]), .QN(n660) );
  DFFRX4 \CNT3_reg[4]  ( .D(n845), .CK(clk), .RN(n1813), .Q(CNT3[4]), .QN(n659) );
  DFFRX4 \CNT3_reg[5]  ( .D(n844), .CK(clk), .RN(n1813), .Q(CNT3[5]), .QN(n658) );
  DFFRX4 \CNT3_reg[6]  ( .D(n843), .CK(clk), .RN(n1813), .Q(CNT3[6]), .QN(n657) );
  DFFRX4 \CNT3_reg[7]  ( .D(n842), .CK(clk), .RN(n1810), .Q(CNT3[7]), .QN(n656) );
  DFFRX4 \CNT1_reg[0]  ( .D(n833), .CK(clk), .RN(n1811), .Q(CNT1[0]), .QN(n647) );
  DFFRX1 \compare_cnt_reg[0]  ( .D(n821), .CK(clk), .RN(n1811), .Q(n3109), 
        .QN(n1738) );
  DFFRX1 compare_all_reg ( .D(n761), .CK(clk), .RN(n1806), .Q(n3077), .QN(
        n1737) );
  DFFRX1 \tree_mem_reg[1]  ( .D(n823), .CK(clk), .RN(n1811), .Q(tree_mem[1]), 
        .QN(n1736) );
  DFFRX1 re_order_en_reg ( .D(n825), .CK(clk), .RN(n1804), .Q(re_order_en), 
        .QN(n1732) );
  DFFRX1 \tree_mem_back_reg[2]  ( .D(n783), .CK(clk), .RN(n1811), .Q(
        tree_mem_back[2]), .QN(n1727) );
  DFFRX1 \state_reg[1]  ( .D(next_state[1]), .CK(clk), .RN(n2914), .Q(state[1]), .QN(n1725) );
  DFFRX1 \com_after_1_reg[0]  ( .D(n811), .CK(clk), .RN(n1809), .Q(
        com_after_1[0]), .QN(n629) );
  DFFRX1 hcode1_1_reg ( .D(n705), .CK(clk), .RN(n1807), .Q(n3061), .QN(n1723)
         );
  DFFRX1 \hcode4_1_reg[0]  ( .D(n723), .CK(clk), .RN(n1805), .Q(n3062), .QN(
        n1721) );
  DFFRX1 \compare_cnt_reg[1]  ( .D(n820), .CK(clk), .RN(n1806), .Q(n3110), 
        .QN(n1720) );
  DFFRX1 \tree_mem_reg[0]  ( .D(n824), .CK(clk), .RN(n1804), .Q(tree_mem[0]), 
        .QN(n1715) );
  DFFRX1 \hcode2_1_reg[1]  ( .D(n772), .CK(clk), .RN(n1811), .Q(n3057), .QN(
        n1713) );
  DFFRX1 \state_reg[0]  ( .D(next_state[0]), .CK(clk), .RN(n1811), .Q(state[0]), .QN(n1712) );
  DFFRX1 \state_reg[2]  ( .D(next_state[2]), .CK(clk), .RN(n1804), .Q(state[2]), .QN(n1711) );
  DFFRX1 \hcode5_1_reg[2]  ( .D(n765), .CK(clk), .RN(n1811), .Q(n3056), .QN(
        n1709) );
  DFFRX1 \hcode5_1_reg[3]  ( .D(n766), .CK(clk), .RN(n1804), .Q(n3053), .QN(
        n1708) );
  DFFRX1 \hcode6_reg[2]  ( .D(n708), .CK(clk), .RN(n1812), .Q(n3066), .QN(
        n1707) );
  DFFRX1 \hcode5_reg[1]  ( .D(n768), .CK(clk), .RN(n1804), .Q(n3070), .QN(
        n1706) );
  DFFRX1 \hcode5_1_reg[1]  ( .D(n764), .CK(clk), .RN(n1804), .Q(n3059), .QN(
        n1705) );
  DFFRX1 \tree_mem_reg[2]  ( .D(n822), .CK(clk), .RN(n2914), .Q(tree_mem[2]), 
        .QN(n1702) );
  DFFRX1 \hcode5_reg[2]  ( .D(n769), .CK(clk), .RN(n1804), .Q(n3067), .QN(
        n1699) );
  DFFRX1 \hcode6_1_reg[2]  ( .D(n758), .CK(clk), .RN(n1807), .Q(n3055), .QN(
        n1698) );
  DFFRX1 \hcode6_1_reg[3]  ( .D(n759), .CK(clk), .RN(n1806), .Q(n3052), .QN(
        n1697) );
  DFFRX1 \hcode6_reg[1]  ( .D(n707), .CK(clk), .RN(n1812), .Q(n3071), .QN(
        n1696) );
  TLATX1 \next_state_reg[1]  ( .G(N202), .D(N204), .Q(next_state[1]) );
  TLATX1 \next_state_reg[2]  ( .G(N202), .D(N205), .Q(next_state[2]) );
  TLATX1 \next_state_reg[0]  ( .G(N202), .D(N203), .Q(next_state[0]) );
  TLATX1 \M1_1_reg[4]  ( .G(N644), .D(N654), .Q(n3103) );
  TLATX1 \M1_1_reg[3]  ( .G(N644), .D(N653), .Q(n3104) );
  TLATX1 \M1_1_reg[2]  ( .G(N644), .D(N652), .Q(n3105) );
  TLATX1 \M1_1_reg[1]  ( .G(N644), .D(N651), .Q(n3106) );
  TLATX1 \M1_1_reg[0]  ( .G(N644), .D(N650), .Q(n3107) );
  TLATX1 \M3_1_reg[4]  ( .G(N672), .D(N682), .Q(n3093) );
  TLATX1 \M3_1_reg[3]  ( .G(N672), .D(N681), .Q(n3094) );
  TLATX1 \M3_1_reg[2]  ( .G(N672), .D(N680), .Q(n3095) );
  TLATX1 \M3_1_reg[1]  ( .G(N672), .D(N679), .Q(n3096) );
  TLATX1 \M3_1_reg[0]  ( .G(N672), .D(N678), .Q(n3097) );
  TLATXL \M6_1_reg[4]  ( .G(N714), .D(N724), .Q(n3078) );
  TLATXL \M6_1_reg[3]  ( .G(N714), .D(N723), .Q(n3079) );
  TLATXL \M6_1_reg[2]  ( .G(N714), .D(N722), .Q(n3080) );
  TLATXL \M6_1_reg[1]  ( .G(N714), .D(N721), .Q(n3081) );
  TLATXL \M6_1_reg[0]  ( .G(N714), .D(N720), .Q(n3082) );
  TLATXL \M2_1_reg[4]  ( .G(N658), .D(N668), .Q(n3098) );
  TLATXL \M2_1_reg[3]  ( .G(N658), .D(N667), .Q(n3099) );
  TLATXL \M2_1_reg[2]  ( .G(N658), .D(N666), .Q(n3100) );
  TLATXL \M2_1_reg[1]  ( .G(N658), .D(N665), .Q(n3101) );
  TLATXL \M2_1_reg[0]  ( .G(N658), .D(N664), .Q(n3102) );
  TLATXL \M5_1_reg[4]  ( .G(N700), .D(N710), .Q(n3083) );
  TLATXL \M5_1_reg[3]  ( .G(N700), .D(N709), .Q(n3084) );
  TLATXL \M5_1_reg[2]  ( .G(N700), .D(N708), .Q(n3085) );
  TLATXL \M5_1_reg[1]  ( .G(N700), .D(N707), .Q(n3086) );
  TLATXL \M5_1_reg[0]  ( .G(N700), .D(N706), .Q(n3087) );
  TLATXL \M4_1_reg[4]  ( .G(N686), .D(N696), .Q(n3088) );
  TLATXL \M4_1_reg[3]  ( .G(N686), .D(N695), .Q(n3089) );
  TLATXL \M4_1_reg[2]  ( .G(N686), .D(N694), .Q(n3090) );
  TLATXL \M4_1_reg[1]  ( .G(N686), .D(N693), .Q(n3091) );
  TLATXL \M4_1_reg[0]  ( .G(N686), .D(N692), .Q(n3092) );
  DFFRX2 \hcode5_reg[0]  ( .D(n770), .CK(clk), .RN(n1804), .Q(n3049), .QN(
        n1704) );
  DFFRX1 out_en_reg ( .D(n762), .CK(clk), .RN(n1807), .Q(out_en) );
  DFFRX1 \hcode6_reg[0]  ( .D(n706), .CK(clk), .RN(n1811), .Q(n3076), .QN(
        n1695) );
  DFFRX1 \hcode6_1_reg[1]  ( .D(n757), .CK(clk), .RN(n1805), .Q(n3060), .QN(
        n1118) );
  DFFRX1 \hcode6_1_reg[4]  ( .D(n760), .CK(clk), .RN(n1805), .QN(n1115) );
  DFFRX1 \hcode5_reg[3]  ( .D(n695), .CK(clk), .RN(n1812), .QN(n1114) );
  DFFRX1 \hcode6_reg[3]  ( .D(n694), .CK(clk), .RN(n1812), .QN(n1097) );
  DFFRX1 \hcode5_reg[4]  ( .D(n691), .CK(clk), .RN(n1812), .QN(n1113) );
  DFFRX1 \hcode6_reg[4]  ( .D(n690), .CK(clk), .RN(n1812), .QN(n1096) );
  DFFRX1 \hcode4_1_reg[3]  ( .D(n738), .CK(clk), .RN(n1812), .Q(n3051) );
  DFFRX1 \hcode4_1_reg[2]  ( .D(n733), .CK(clk), .RN(n1812), .Q(n3054) );
  DFFRX1 \hcode4_1_reg[1]  ( .D(n728), .CK(clk), .RN(n1807), .Q(n3058) );
  DFFRX1 \hcode2_reg[1]  ( .D(n696), .CK(clk), .RN(n1812), .Q(n3068), .QN(
        n1733) );
  DFFRX1 \hcode2_1_reg[0]  ( .D(n771), .CK(clk), .RN(n1804), .QN(n1731) );
  DFFRX1 \hcode3_1_reg[1]  ( .D(n779), .CK(clk), .RN(n1804), .QN(n1722) );
  DFFRX1 \hcode3_1_reg[3]  ( .D(n781), .CK(clk), .RN(n2914), .QN(n1718) );
  DFFRX1 \hcode3_reg[2]  ( .D(n693), .CK(clk), .RN(n1812), .Q(n3065), .QN(
        n1717) );
  DFFRX1 \hcode3_1_reg[2]  ( .D(n780), .CK(clk), .RN(n1806), .QN(n1716) );
  DFFRX1 \hcode3_1_reg[0]  ( .D(n778), .CK(clk), .RN(n1811), .QN(n1730) );
  DFFRX1 \hcode6_1_reg[0]  ( .D(n756), .CK(clk), .RN(n1806), .Q(n3063), .QN(
        n1701) );
  DFFRX1 \hcode4_reg[1]  ( .D(n777), .CK(clk), .RN(n1813), .Q(n3069), .QN(
        n1739) );
  DFFRX1 \hcode5_1_reg[0]  ( .D(n763), .CK(clk), .RN(n1804), .Q(n3050), .QN(
        n1693) );
  DFFRX1 \hcode5_1_reg[4]  ( .D(n767), .CK(clk), .RN(n1811), .QN(n1703) );
  DFFRX1 \com_after_1_reg[6]  ( .D(n817), .CK(clk), .RN(n1808), .Q(
        com_after_1[6]), .QN(n635) );
  DFFRX1 \com_after_1_reg[3]  ( .D(n814), .CK(clk), .RN(n1808), .Q(
        com_after_1[3]), .QN(n632) );
  DFFRX1 \com_after_1_reg[4]  ( .D(n815), .CK(clk), .RN(n1809), .Q(
        com_after_1[4]), .QN(n633) );
  DFFRX1 \com_after_1_reg[5]  ( .D(n816), .CK(clk), .RN(n1808), .Q(
        com_after_1[5]), .QN(n634) );
  DFFRX1 \tree_mem_back_reg[0]  ( .D(n785), .CK(clk), .RN(n1804), .Q(
        tree_mem_back[0]), .QN(n1734) );
  DFFRX2 \CNT4_reg[0]  ( .D(n865), .CK(clk), .RN(n1804), .Q(CNT4[0]), .QN(n679) );
  DFFRX4 \CNT5_reg[5]  ( .D(n852), .CK(clk), .RN(n1810), .Q(CNT5[5]), .QN(n666) );
  DFFRX4 \CNT5_reg[4]  ( .D(n853), .CK(clk), .RN(n1810), .Q(CNT5[4]), .QN(n667) );
  DFFRX4 \CNT5_reg[3]  ( .D(n854), .CK(clk), .RN(n1810), .Q(CNT5[3]), .QN(n668) );
  DFFRX4 \CNT6_reg[4]  ( .D(n869), .CK(clk), .RN(n1810), .Q(CNT6[4]), .QN(n683) );
  DFFRX2 \CNT5_reg[2]  ( .D(n855), .CK(clk), .RN(n1810), .Q(CNT5[2]), .QN(n669) );
  DFFRX4 \CNT6_reg[7]  ( .D(n866), .CK(clk), .RN(n1809), .Q(CNT6[7]), .QN(n680) );
  DFFRX2 \CNT6_reg[5]  ( .D(n868), .CK(clk), .RN(n1809), .Q(CNT6[5]), .QN(n682) );
  DFFRX2 \CNT6_reg[3]  ( .D(n870), .CK(clk), .RN(n1808), .Q(CNT6[3]), .QN(n684) );
  DFFRX2 \CNT6_reg[6]  ( .D(n867), .CK(clk), .RN(n1810), .Q(CNT6[6]), .QN(n681) );
  DFFRX2 \tree_mem_back_reg[1]  ( .D(n784), .CK(clk), .RN(n1805), .Q(
        tree_mem_back[1]), .QN(n1741) );
  DFFRX2 \CNT6_reg[2]  ( .D(n871), .CK(clk), .RN(n1809), .Q(CNT6[2]), .QN(n685) );
  DFFRX2 \CNT5_reg[6]  ( .D(n851), .CK(clk), .RN(n1810), .Q(CNT5[6]), .QN(n665) );
  TLATX2 \HC1_reg[1]  ( .G(N644), .D(N646), .Q(HC1[1]) );
  TLATX2 \HC1_reg[2]  ( .G(N644), .D(N647), .Q(HC1[2]) );
  TLATX2 \HC1_reg[3]  ( .G(N644), .D(N648), .Q(HC1[3]) );
  TLATX2 \HC1_reg[4]  ( .G(N644), .D(N649), .Q(HC1[4]) );
  TLATX2 \HC1_reg[0]  ( .G(N644), .D(N645), .Q(HC1[0]) );
  TLATX2 \HC5_reg[1]  ( .G(N700), .D(N702), .Q(HC5[1]) );
  TLATX2 \HC5_reg[2]  ( .G(N700), .D(N703), .Q(HC5[2]) );
  TLATX2 \HC5_reg[3]  ( .G(N700), .D(N704), .Q(HC5[3]) );
  TLATX2 \HC5_reg[4]  ( .G(N700), .D(N705), .Q(HC5[4]) );
  TLATX2 \HC5_reg[0]  ( .G(N700), .D(N701), .Q(HC5[0]) );
  DFFRX2 \hcode4_reg[3]  ( .D(n692), .CK(clk), .RN(n1812), .QN(n1694) );
  DFFRX2 \CNT6_reg[1]  ( .D(n872), .CK(clk), .RN(n1810), .Q(CNT6[1]), .QN(n686) );
  DFFRX2 \CNT6_reg[0]  ( .D(n873), .CK(clk), .RN(n1810), .Q(CNT6[0]), .QN(n687) );
  DFFRX2 \CNT5_reg[0]  ( .D(n857), .CK(clk), .RN(n1809), .Q(CNT5[0]), .QN(n671) );
  DFFRX4 \CNT5_reg[7]  ( .D(n850), .CK(clk), .RN(n1809), .Q(CNT5[7]), .QN(n664) );
  DFFRX2 \com_after_1_reg[1]  ( .D(n812), .CK(clk), .RN(n1809), .Q(
        com_after_1[1]), .QN(n630) );
  TLATXL \HC4_reg[1]  ( .G(N686), .D(N688), .QN(n1126) );
  TLATXL \HC4_reg[2]  ( .G(N686), .D(N689), .QN(n1127) );
  TLATXL \HC4_reg[3]  ( .G(N686), .D(N690), .QN(n1128) );
  TLATXL \HC4_reg[4]  ( .G(N686), .D(N691), .QN(n1129) );
  TLATXL \HC4_reg[0]  ( .G(N686), .D(N687), .QN(n1125) );
  TLATXL \HC6_reg[1]  ( .G(N714), .D(N716), .QN(n1122) );
  TLATXL \HC2_reg[1]  ( .G(N658), .D(N660), .QN(n1131) );
  TLATX2 \HC6_reg[2]  ( .G(N714), .D(N717), .Q(HC6[2]) );
  TLATX2 \HC2_reg[2]  ( .G(N658), .D(N661), .Q(HC2[2]) );
  TLATXL \HC6_reg[3]  ( .G(N714), .D(N718), .QN(n1123) );
  TLATXL \HC2_reg[3]  ( .G(N658), .D(N662), .QN(n1132) );
  TLATXL \HC6_reg[4]  ( .G(N714), .D(N719), .QN(n1124) );
  TLATXL \HC2_reg[4]  ( .G(N658), .D(N663), .QN(n1133) );
  TLATXL \HC6_reg[0]  ( .G(N714), .D(N715), .QN(n1121) );
  TLATXL \HC2_reg[0]  ( .G(N658), .D(N659), .QN(n1130) );
  TLATX2 \HC3_reg[1]  ( .G(N672), .D(N674), .Q(HC3[1]) );
  TLATX2 \HC3_reg[2]  ( .G(N672), .D(N675), .Q(HC3[2]) );
  TLATX2 \HC3_reg[3]  ( .G(N672), .D(N676), .Q(HC3[3]) );
  TLATX2 \HC3_reg[4]  ( .G(N672), .D(N677), .Q(HC3[4]) );
  TLATX2 \HC3_reg[0]  ( .G(N672), .D(N673), .Q(HC3[0]) );
  DFFRX2 CNT_valid_reg ( .D(n755), .CK(clk), .RN(n1807), .Q(CNT_valid), .QN(
        n579) );
  DFFRX2 \M6_reg[4]  ( .D(n742), .CK(clk), .RN(n1807), .Q(M6[4]), .QN(n553) );
  DFFRX2 \M5_reg[4]  ( .D(n741), .CK(clk), .RN(n1805), .Q(M5[4]), .QN(n551) );
  DFFRX2 \M3_reg[4]  ( .D(n740), .CK(clk), .RN(n1805), .Q(M3[4]), .QN(n549) );
  DFFRX2 \M2_reg[4]  ( .D(n739), .CK(clk), .RN(n1805), .Q(M2[4]), .QN(n547) );
  DFFRX2 \M6_reg[3]  ( .D(n737), .CK(clk), .RN(n1812), .Q(M6[3]), .QN(n544) );
  DFFRX2 \M5_reg[3]  ( .D(n736), .CK(clk), .RN(n1812), .Q(M5[3]), .QN(n542) );
  DFFRX2 \M3_reg[3]  ( .D(n735), .CK(clk), .RN(n1812), .Q(M3[3]), .QN(n540) );
  DFFRX2 \M2_reg[3]  ( .D(n734), .CK(clk), .RN(n1807), .Q(M2[3]), .QN(n538) );
  DFFRX2 \M6_reg[2]  ( .D(n732), .CK(clk), .RN(n1807), .Q(M6[2]), .QN(n535) );
  DFFRX2 \M5_reg[2]  ( .D(n731), .CK(clk), .RN(n1812), .Q(M5[2]), .QN(n533) );
  DFFRX2 \M3_reg[2]  ( .D(n730), .CK(clk), .RN(n1807), .Q(M3[2]), .QN(n531) );
  DFFRX2 \M2_reg[2]  ( .D(n729), .CK(clk), .RN(n1807), .Q(M2[2]), .QN(n529) );
  DFFRX2 \M6_reg[1]  ( .D(n727), .CK(clk), .RN(n1807), .Q(M6[1]), .QN(n526) );
  DFFRX2 \M5_reg[1]  ( .D(n726), .CK(clk), .RN(n1805), .Q(M5[1]), .QN(n524) );
  DFFRX2 \M3_reg[1]  ( .D(n725), .CK(clk), .RN(n1805), .Q(M3[1]), .QN(n522) );
  DFFRX2 \M2_reg[1]  ( .D(n724), .CK(clk), .RN(n1805), .Q(M2[1]), .QN(n520) );
  DFFRX2 \M4_reg[4]  ( .D(n719), .CK(clk), .RN(n1806), .Q(M4[4]), .QN(n511) );
  DFFRX2 \M4_reg[3]  ( .D(n718), .CK(clk), .RN(n1806), .Q(M4[3]), .QN(n509) );
  DFFRX2 \M4_reg[2]  ( .D(n717), .CK(clk), .RN(n1806), .Q(M4[2]), .QN(n507) );
  DFFRX2 \M4_reg[1]  ( .D(n716), .CK(clk), .RN(n1806), .Q(M4[1]), .QN(n505) );
  DFFRX2 \M1_reg[4]  ( .D(n712), .CK(clk), .RN(n1812), .Q(M1[4]), .QN(n497) );
  DFFRX2 \M1_reg[3]  ( .D(n711), .CK(clk), .RN(n1812), .Q(M1[3]), .QN(n495) );
  DFFRX2 \M1_reg[2]  ( .D(n710), .CK(clk), .RN(n1812), .Q(M1[2]), .QN(n493) );
  DFFRX2 \M1_reg[1]  ( .D(n709), .CK(clk), .RN(n1812), .Q(M1[1]), .QN(n491) );
  DFFRX2 \M6_reg[0]  ( .D(n704), .CK(clk), .RN(n1812), .Q(M6[0]), .QN(n485) );
  DFFRX2 \M5_reg[0]  ( .D(n703), .CK(clk), .RN(n1812), .Q(M5[0]), .QN(n483) );
  DFFRX2 \M4_reg[0]  ( .D(n702), .CK(clk), .RN(n1812), .Q(M4[0]), .QN(n481) );
  DFFRX2 \M3_reg[0]  ( .D(n701), .CK(clk), .RN(n1812), .Q(M3[0]), .QN(n479) );
  DFFRX2 \M2_reg[0]  ( .D(n700), .CK(clk), .RN(n1812), .Q(M2[0]), .QN(n477) );
  DFFRX2 \M1_reg[0]  ( .D(n699), .CK(clk), .RN(n1812), .Q(M1[0]), .QN(n475) );
  DFFRX2 code_valid_reg ( .D(n698), .CK(clk), .RN(n1812), .Q(code_valid), .QN(
        n474) );
  DFFRX2 \com_after_1_reg[2]  ( .D(n813), .CK(clk), .RN(n1809), .Q(
        com_after_1[2]), .QN(n631) );
  DFFRHQX8 \CNT1_reg[1]  ( .D(n832), .CK(clk), .RN(n1807), .Q(n1243) );
  DFFRHQX8 \CNT1_reg[3]  ( .D(n830), .CK(clk), .RN(n1811), .Q(n1242) );
  DFFRHQX8 \CNT2_reg[1]  ( .D(n840), .CK(clk), .RN(n1813), .Q(n1241) );
  DFFRHQX8 \CNT2_reg[7]  ( .D(n834), .CK(clk), .RN(n1813), .Q(n1238) );
  DFFRHQX8 \CNT2_reg[6]  ( .D(n835), .CK(clk), .RN(n1808), .Q(n1236) );
  DFFRHQX8 \CNT2_reg[3]  ( .D(n838), .CK(clk), .RN(n1813), .Q(n1235) );
  DFFRHQX8 \CNT1_reg[7]  ( .D(n826), .CK(clk), .RN(n1808), .Q(n1229) );
  DFFRHQX8 \CNT1_reg[5]  ( .D(n828), .CK(clk), .RN(n1811), .Q(n1227) );
  DFFRHQX8 \CNT2_reg[0]  ( .D(n841), .CK(clk), .RN(n1808), .Q(n1213) );
  DFFRHQX8 \CNT2_reg[2]  ( .D(n839), .CK(clk), .RN(n1808), .Q(n1212) );
  DFFRHQX8 \CNT2_reg[4]  ( .D(n837), .CK(clk), .RN(n1808), .Q(n1210) );
  DFFRHQX8 \CNT2_reg[5]  ( .D(n836), .CK(clk), .RN(n1808), .Q(n1207) );
  DFFRHQX8 \CNT1_reg[2]  ( .D(n831), .CK(clk), .RN(n1809), .Q(n1206) );
  DFFRHQX8 \CNT1_reg[4]  ( .D(n829), .CK(clk), .RN(n1811), .Q(n1204) );
  DFFRX2 \CNT3_reg[0]  ( .D(n849), .CK(clk), .RN(n1810), .Q(CNT3[0]), .QN(n663) );
  DFFRX2 \CNT4_reg[1]  ( .D(n864), .CK(clk), .RN(n1804), .Q(CNT4[1]), .QN(n678) );
  DFFRX2 \CNT4_reg[6]  ( .D(n859), .CK(clk), .RN(n1805), .Q(CNT4[6]), .QN(n673) );
  DFFRX4 \CNT4_reg[5]  ( .D(n860), .CK(clk), .RN(n1809), .Q(CNT4[5]), .QN(n674) );
  DFFRHQX4 \CNT1_reg[6]  ( .D(n827), .CK(clk), .RN(n1811), .Q(n1244) );
  DFFRX2 \CNT5_reg[1]  ( .D(n856), .CK(clk), .RN(n1810), .Q(CNT5[1]), .QN(n670) );
  NOR2X4 U1037 ( .A(n942), .B(n2237), .Y(n936) );
  NAND3X6 U1038 ( .A(n943), .B(n940), .C(n936), .Y(n934) );
  BUFX20 U1039 ( .A(n933), .Y(n930) );
  NAND2X8 U1040 ( .A(n932), .B(n931), .Y(n933) );
  NAND2X6 U1041 ( .A(n934), .B(n938), .Y(n931) );
  NAND2X6 U1042 ( .A(n935), .B(n1111), .Y(n932) );
  MXI2X4 U1043 ( .A(n1322), .B(n1192), .S0(n930), .Y(n2613) );
  NAND3X6 U1044 ( .A(n943), .B(n941), .C(n940), .Y(n935) );
  NAND3X8 U1045 ( .A(n2241), .B(n2240), .C(n2239), .Y(n940) );
  NOR2X8 U1046 ( .A(n2238), .B(n1779), .Y(n942) );
  NAND3X8 U1047 ( .A(n1710), .B(n2220), .C(n2221), .Y(n943) );
  CLKINVX20 U1048 ( .A(n937), .Y(n1796) );
  BUFX8 U1049 ( .A(n1795), .Y(n937) );
  CLKINVX8 U1050 ( .A(n939), .Y(n938) );
  NAND2X6 U1051 ( .A(n2243), .B(n2422), .Y(n939) );
  MXI2X4 U1052 ( .A(n2398), .B(n2397), .S0(n1795), .Y(n2422) );
  NOR2X6 U1053 ( .A(n942), .B(n2228), .Y(n941) );
  INVX3 U1054 ( .A(n1633), .Y(n1632) );
  NOR2X4 U1055 ( .A(n1043), .B(n1041), .Y(n1033) );
  NOR2X4 U1056 ( .A(n1043), .B(n1042), .Y(n1036) );
  CLKINVX20 U1057 ( .A(n1023), .Y(n1790) );
  NOR2X4 U1058 ( .A(n948), .B(n944), .Y(n2186) );
  NOR2X2 U1059 ( .A(n1761), .B(n2190), .Y(n944) );
  BUFX4 U1060 ( .A(n2179), .Y(n945) );
  NAND2X8 U1061 ( .A(n1032), .B(n1039), .Y(n1031) );
  NAND2X8 U1062 ( .A(n2072), .B(n1431), .Y(n1477) );
  AND2X6 U1063 ( .A(n2033), .B(n2034), .Y(n1685) );
  INVX4 U1064 ( .A(n2592), .Y(n2594) );
  NOR2X8 U1065 ( .A(n1650), .B(n946), .Y(n1555) );
  NOR2X8 U1066 ( .A(n1775), .B(n1389), .Y(n946) );
  BUFX4 U1067 ( .A(n2184), .Y(n947) );
  NOR2X2 U1068 ( .A(n2295), .B(n2208), .Y(n948) );
  NAND2X4 U1069 ( .A(n2174), .B(n2265), .Y(n2149) );
  BUFX4 U1070 ( .A(n2164), .Y(n949) );
  INVX12 U1071 ( .A(n2179), .Y(n2085) );
  BUFX4 U1072 ( .A(n2171), .Y(n950) );
  BUFX4 U1073 ( .A(n1224), .Y(n951) );
  NOR2X8 U1074 ( .A(n1990), .B(n1405), .Y(n1043) );
  CLKINVX12 U1075 ( .A(n958), .Y(n1195) );
  INVX6 U1076 ( .A(n2076), .Y(n1551) );
  INVX12 U1077 ( .A(n952), .Y(n1989) );
  CLKAND2X8 U1078 ( .A(n2093), .B(n1980), .Y(n952) );
  BUFX4 U1079 ( .A(n2266), .Y(n953) );
  BUFX4 U1080 ( .A(n2254), .Y(n954) );
  INVX8 U1081 ( .A(n1290), .Y(n2059) );
  NAND2X4 U1082 ( .A(n1302), .B(n1649), .Y(n958) );
  INVX12 U1083 ( .A(n1022), .Y(n2254) );
  BUFX4 U1084 ( .A(n2173), .Y(n955) );
  NAND2X8 U1085 ( .A(n2171), .B(n2172), .Y(n1274) );
  NOR2X6 U1086 ( .A(n970), .B(n956), .Y(n969) );
  OAI21X4 U1087 ( .A0(n2059), .A1(n1764), .B0(n2050), .Y(n956) );
  INVX8 U1088 ( .A(n1473), .Y(n1774) );
  BUFX4 U1089 ( .A(n1970), .Y(n957) );
  NAND4X8 U1090 ( .A(n1554), .B(n1549), .C(n1248), .D(n1628), .Y(n1552) );
  NAND2X8 U1091 ( .A(n1385), .B(n1387), .Y(n1474) );
  NOR2X8 U1092 ( .A(n1386), .B(n1079), .Y(n1385) );
  OAI2BB1X4 U1093 ( .A0N(n1760), .A1N(n2092), .B0(n1059), .Y(n1068) );
  BUFX20 U1094 ( .A(n1786), .Y(n1356) );
  MXI2X6 U1095 ( .A(n678), .B(n1064), .S0(n1356), .Y(n1954) );
  BUFX16 U1096 ( .A(n2576), .Y(n1383) );
  NAND3X8 U1097 ( .A(n1554), .B(n1550), .C(n1549), .Y(n1548) );
  BUFX4 U1098 ( .A(n1984), .Y(n959) );
  AND2X8 U1099 ( .A(n1081), .B(n1396), .Y(n1619) );
  MXI2X4 U1100 ( .A(n961), .B(n960), .S0(n1790), .Y(n1396) );
  CLKINVX6 U1101 ( .A(n2074), .Y(n960) );
  CLKINVX6 U1102 ( .A(n2073), .Y(n961) );
  NAND3X6 U1103 ( .A(n1037), .B(n1038), .C(n1033), .Y(n1032) );
  NAND2X6 U1104 ( .A(n1427), .B(n1426), .Y(n987) );
  NAND2X6 U1105 ( .A(n1936), .B(n1103), .Y(n1656) );
  INVX3 U1106 ( .A(n1919), .Y(n1920) );
  INVX8 U1107 ( .A(n2009), .Y(n1332) );
  MXI2X4 U1108 ( .A(n963), .B(n962), .S0(n1024), .Y(n2009) );
  CLKINVX6 U1109 ( .A(n1026), .Y(n962) );
  CLKINVX6 U1110 ( .A(n1913), .Y(n963) );
  MXI2X2 U1111 ( .A(CNT2[2]), .B(CNT1[2]), .S0(n1343), .Y(n1934) );
  NAND2X8 U1112 ( .A(n1001), .B(n1931), .Y(n1017) );
  NAND2X6 U1113 ( .A(n1675), .B(n1017), .Y(n1598) );
  OR2X8 U1114 ( .A(n1980), .B(n2093), .Y(n1303) );
  NOR2X8 U1115 ( .A(n1591), .B(n1590), .Y(n1622) );
  BUFX4 U1116 ( .A(n1952), .Y(n964) );
  INVX12 U1117 ( .A(n1073), .Y(n1771) );
  AND2X8 U1118 ( .A(n2064), .B(n1419), .Y(n1194) );
  BUFX4 U1119 ( .A(n1016), .Y(n965) );
  NAND2X8 U1120 ( .A(n2158), .B(n2157), .Y(n1430) );
  AND2X8 U1121 ( .A(n2181), .B(n2259), .Y(n1644) );
  INVX8 U1122 ( .A(n2078), .Y(n1547) );
  AND2X8 U1123 ( .A(n1366), .B(n1311), .Y(n1365) );
  NAND3X6 U1124 ( .A(n1295), .B(n1090), .C(n1603), .Y(n1599) );
  NAND3X8 U1125 ( .A(n1327), .B(n966), .C(n1516), .Y(n1940) );
  NOR2X8 U1126 ( .A(n1511), .B(n1513), .Y(n966) );
  INVX12 U1127 ( .A(n1917), .Y(n967) );
  NAND2X4 U1128 ( .A(n967), .B(n675), .Y(n1434) );
  INVX16 U1129 ( .A(n1517), .Y(n1952) );
  CLKBUFX3 U1130 ( .A(n1967), .Y(n968) );
  NAND3X4 U1131 ( .A(n1280), .B(n951), .C(n2045), .Y(n1676) );
  NAND3X6 U1132 ( .A(n1678), .B(n1677), .C(n1676), .Y(n2248) );
  NAND3X8 U1133 ( .A(n1372), .B(n969), .C(n1371), .Y(n1380) );
  NOR2X4 U1134 ( .A(n2134), .B(n2055), .Y(n970) );
  NAND3X6 U1135 ( .A(n2121), .B(n2122), .C(CNT6[7]), .Y(n1531) );
  BUFX20 U1136 ( .A(n1646), .Y(n1673) );
  BUFX12 U1137 ( .A(n1646), .Y(n1374) );
  NAND2X8 U1138 ( .A(n971), .B(n2075), .Y(n1633) );
  NAND2X8 U1139 ( .A(n1619), .B(n2077), .Y(n971) );
  NAND3X8 U1140 ( .A(n2022), .B(n2021), .C(CNT5[7]), .Y(n2023) );
  BUFX4 U1141 ( .A(n1367), .Y(n972) );
  BUFX4 U1142 ( .A(n1915), .Y(n973) );
  BUFX4 U1143 ( .A(n1673), .Y(n974) );
  NAND2X6 U1144 ( .A(n2162), .B(n953), .Y(n1498) );
  BUFX4 U1145 ( .A(n2392), .Y(n975) );
  CLKBUFX12 U1146 ( .A(n1803), .Y(n1352) );
  NOR2X8 U1147 ( .A(n1668), .B(n1166), .Y(n1162) );
  BUFX4 U1148 ( .A(\com[4][3] ), .Y(n976) );
  CLKBUFX20 U1149 ( .A(n1801), .Y(n979) );
  NAND2X2 U1150 ( .A(n979), .B(n2393), .Y(n1522) );
  MXI2X8 U1151 ( .A(n1192), .B(n1322), .S0(n1313), .Y(\com[3][4] ) );
  CLKBUFX16 U1152 ( .A(n1801), .Y(n1313) );
  BUFX16 U1153 ( .A(n933), .Y(n1801) );
  MXI2X6 U1154 ( .A(n2400), .B(n2399), .S0(n1796), .Y(n2614) );
  BUFX4 U1155 ( .A(n2413), .Y(n977) );
  BUFX4 U1156 ( .A(n2386), .Y(n978) );
  INVX6 U1157 ( .A(n2596), .Y(n2450) );
  BUFX20 U1158 ( .A(n1785), .Y(n1024) );
  BUFX4 U1159 ( .A(n2057), .Y(n980) );
  BUFX4 U1160 ( .A(n1673), .Y(n981) );
  NAND4X6 U1161 ( .A(n2186), .B(n1061), .C(n2187), .D(n1778), .Y(n986) );
  BUFX20 U1162 ( .A(n1422), .Y(n982) );
  NAND4X8 U1163 ( .A(n987), .B(n986), .C(n984), .D(n983), .Y(n1422) );
  NAND2X8 U1164 ( .A(n1424), .B(n1563), .Y(n983) );
  NAND2X8 U1165 ( .A(n1423), .B(n985), .Y(n984) );
  CLKINVX6 U1166 ( .A(n1661), .Y(n985) );
  MXI2X4 U1167 ( .A(n2202), .B(n2292), .S0(n982), .Y(n2388) );
  AND2X8 U1168 ( .A(n2155), .B(n2154), .Y(n1060) );
  AND2X6 U1169 ( .A(n2434), .B(n990), .Y(n1670) );
  MXI2X8 U1170 ( .A(n992), .B(n991), .S0(n930), .Y(n2434) );
  CLKINVX20 U1171 ( .A(n2611), .Y(n988) );
  DLY3X1 U1172 ( .A(n2434), .Y(n989) );
  INVX6 U1173 ( .A(n2611), .Y(n990) );
  OR2X8 U1174 ( .A(n2434), .B(n988), .Y(n2428) );
  CLKINVX4 U1175 ( .A(n978), .Y(n991) );
  INVX12 U1176 ( .A(n1283), .Y(n992) );
  CLKAND2X12 U1177 ( .A(n2301), .B(n2302), .Y(n1187) );
  NAND3X2 U1178 ( .A(n2300), .B(n632), .C(\com[3][3] ), .Y(n2301) );
  NAND2X8 U1179 ( .A(n2303), .B(n1187), .Y(n1186) );
  NAND2X8 U1180 ( .A(n1009), .B(n2036), .Y(n1074) );
  NAND2X8 U1181 ( .A(n2035), .B(n1685), .Y(n2036) );
  INVXL U1183 ( .A(n979), .Y(n994) );
  CLKINVX1 U1184 ( .A(n994), .Y(n995) );
  NAND2X2 U1187 ( .A(n1801), .B(n1102), .Y(n2401) );
  NOR2X8 U1190 ( .A(n1464), .B(n607), .Y(n2631) );
  NAND2X6 U1192 ( .A(n1053), .B(n791), .Y(n1453) );
  INVX4 U1193 ( .A(n2300), .Y(n1320) );
  OR2X6 U1194 ( .A(\com[3][4] ), .B(n633), .Y(n2300) );
  INVXL U1196 ( .A(n1352), .Y(n997) );
  CLKINVX1 U1197 ( .A(n997), .Y(n998) );
  NAND2X2 U1199 ( .A(n1352), .B(n2597), .Y(n1411) );
  NOR2X4 U1200 ( .A(n1352), .B(n1412), .Y(n1055) );
  INVX8 U1201 ( .A(n2208), .Y(n2296) );
  INVX8 U1202 ( .A(n2404), .Y(n999) );
  CLKINVX8 U1203 ( .A(n2275), .Y(n2404) );
  OAI22X1 U1206 ( .A0(n2361), .A1(\com[2][5] ), .B0(n2372), .B1(\com[2][4] ), 
        .Y(n2362) );
  AOI2BB2X4 U1207 ( .B0(\com[2][5] ), .B1(n2361), .A0N(n2363), .A1N(n2362), 
        .Y(n1451) );
  INVX1 U1208 ( .A(\com[3][5] ), .Y(n2361) );
  BUFX3 U1210 ( .A(n1978), .Y(n1000) );
  NAND2X8 U1211 ( .A(n1611), .B(n1433), .Y(n1315) );
  NOR2X6 U1212 ( .A(n1089), .B(n1525), .Y(n1276) );
  NAND2X8 U1213 ( .A(n1963), .B(n1964), .Y(n1005) );
  MXI2X4 U1214 ( .A(CNT3[5]), .B(n1928), .S0(n1025), .Y(n1001) );
  MXI2X4 U1215 ( .A(CNT3[5]), .B(n1928), .S0(n1025), .Y(n1975) );
  INVX16 U1216 ( .A(n1360), .Y(n1367) );
  NAND2X8 U1217 ( .A(n2020), .B(n1684), .Y(n2037) );
  BUFX16 U1218 ( .A(n1479), .Y(n1002) );
  AND2X8 U1219 ( .A(n2117), .B(n1082), .Y(n1106) );
  CLKAND2X12 U1220 ( .A(n2117), .B(n1631), .Y(n2125) );
  CLKINVX8 U1221 ( .A(n1089), .Y(n2044) );
  MX2X4 U1222 ( .A(n679), .B(n2007), .S0(n1279), .Y(n1965) );
  OR2X8 U1223 ( .A(n1954), .B(n2052), .Y(n1682) );
  INVX8 U1224 ( .A(n2184), .Y(n1003) );
  INVX12 U1225 ( .A(n2092), .Y(n2184) );
  NAND2X8 U1226 ( .A(n1626), .B(n1553), .Y(n1549) );
  CLKMX2X2 U1227 ( .A(n678), .B(n1064), .S0(n1279), .Y(n1004) );
  CLKINVX1 U1228 ( .A(n2513), .Y(n1006) );
  NOR2X8 U1229 ( .A(n1775), .B(n1389), .Y(n1079) );
  INVXL U1230 ( .A(n1648), .Y(n1007) );
  CLKINVX1 U1231 ( .A(n1007), .Y(n1008) );
  INVX8 U1232 ( .A(n2267), .Y(n2162) );
  CLKINVX3 U1233 ( .A(n2047), .Y(n1399) );
  MXI2XL U1234 ( .A(n2519), .B(n2518), .S0(n1008), .Y(n2522) );
  MXI2XL U1235 ( .A(n2548), .B(n2547), .S0(n1008), .Y(n2667) );
  MXI2XL U1236 ( .A(n2492), .B(n2491), .S0(n1008), .Y(n2509) );
  MXI2XL U1237 ( .A(n2521), .B(n2520), .S0(n1008), .Y(n2575) );
  CLKMX2X3 U1238 ( .A(n661), .B(n1929), .S0(n1025), .Y(n1065) );
  NAND2X8 U1239 ( .A(n1479), .B(n2048), .Y(n1959) );
  NAND3X4 U1240 ( .A(n1989), .B(n1176), .C(n1994), .Y(n1041) );
  NAND3X8 U1241 ( .A(n1575), .B(n1577), .C(n1647), .Y(n2157) );
  NAND2X4 U1242 ( .A(n1583), .B(n1584), .Y(n1273) );
  NAND2X8 U1243 ( .A(n2020), .B(n1684), .Y(n1009) );
  BUFX16 U1244 ( .A(n965), .Y(n1014) );
  NAND2X2 U1245 ( .A(n2118), .B(n685), .Y(n2119) );
  INVX3 U1246 ( .A(n1523), .Y(n1010) );
  INVXL U1247 ( .A(n995), .Y(n1011) );
  CLKINVX1 U1248 ( .A(n1011), .Y(n1012) );
  INVX3 U1249 ( .A(n2140), .Y(n1013) );
  INVX12 U1250 ( .A(n2070), .Y(n2140) );
  INVX4 U1251 ( .A(n2074), .Y(n1062) );
  CLKAND2X12 U1252 ( .A(n2074), .B(n2143), .Y(n2067) );
  INVX8 U1253 ( .A(n2142), .Y(n2074) );
  AND2X8 U1254 ( .A(n1338), .B(CNT6[5]), .Y(n2123) );
  BUFX20 U1255 ( .A(n1217), .Y(n1339) );
  CLKMX2X6 U1256 ( .A(n2113), .B(CNT5[4]), .S0(n1690), .Y(n1391) );
  BUFX2 U1257 ( .A(n1969), .Y(n1018) );
  CLKMX2X6 U1258 ( .A(CNT4[4]), .B(n2003), .S0(n1279), .Y(n1089) );
  NAND2X6 U1259 ( .A(n1172), .B(n1892), .Y(n1895) );
  MXI2X8 U1260 ( .A(n2451), .B(n1147), .S0(n1802), .Y(\com[4][3] ) );
  NAND2X6 U1261 ( .A(n2428), .B(n1409), .Y(n1143) );
  CLKINVX12 U1262 ( .A(n1353), .Y(n1217) );
  NAND3X6 U1263 ( .A(n2027), .B(n2026), .C(n1226), .Y(n2028) );
  NAND3X6 U1264 ( .A(n2027), .B(n1226), .C(n2026), .Y(n2018) );
  INVX8 U1265 ( .A(n2147), .Y(n1015) );
  INVX12 U1266 ( .A(n2257), .Y(n2147) );
  NAND2X2 U1267 ( .A(n2216), .B(n2388), .Y(n2206) );
  INVX6 U1268 ( .A(n2388), .Y(n2217) );
  MX2X6 U1269 ( .A(n1027), .B(n2072), .S0(n1790), .Y(n1016) );
  CLKINVX12 U1270 ( .A(n1790), .Y(n1791) );
  CLKAND2X12 U1271 ( .A(n2038), .B(n2039), .Y(n1997) );
  AND2X8 U1272 ( .A(n1961), .B(n2038), .Y(n1683) );
  NOR2X8 U1273 ( .A(n1961), .B(n2038), .Y(n1266) );
  INVX12 U1274 ( .A(n2038), .Y(n1951) );
  NAND2X6 U1275 ( .A(n2057), .B(n1981), .Y(n1957) );
  INVX8 U1276 ( .A(n1758), .Y(n1479) );
  OAI21X4 U1277 ( .A0(n1937), .A1(n1513), .B0(n1017), .Y(n1608) );
  OR2X8 U1278 ( .A(n1969), .B(n1019), .Y(n1070) );
  CLKINVX6 U1279 ( .A(n1514), .Y(n1019) );
  MXI2X4 U1280 ( .A(n1018), .B(n1020), .S0(n1339), .Y(n1985) );
  CLKINVX6 U1281 ( .A(n1933), .Y(n1020) );
  INVX20 U1282 ( .A(n1021), .Y(n1360) );
  NAND2X8 U1283 ( .A(n1005), .B(n1962), .Y(n1021) );
  INVX4 U1284 ( .A(n1030), .Y(n1431) );
  MXI2X4 U1285 ( .A(n1029), .B(n1028), .S0(n1360), .Y(n1030) );
  NAND2X8 U1286 ( .A(n1302), .B(n1649), .Y(n1023) );
  NAND2X8 U1287 ( .A(n1368), .B(n1417), .Y(n1649) );
  NAND2X8 U1288 ( .A(n1376), .B(n1375), .Y(n1302) );
  CLKMX2X6 U1289 ( .A(n1062), .B(n2143), .S0(n1790), .Y(n1022) );
  BUFX20 U1290 ( .A(n1785), .Y(n1025) );
  NAND2X4 U1291 ( .A(n1332), .B(CNT4[2]), .Y(n1914) );
  CLKINVX6 U1292 ( .A(n1044), .Y(n1026) );
  NAND2X8 U1293 ( .A(n1771), .B(n1030), .Y(n1310) );
  CLKBUFX8 U1294 ( .A(n1030), .Y(n1027) );
  CLKINVX6 U1295 ( .A(n1399), .Y(n1028) );
  CLKINVX6 U1296 ( .A(n1398), .Y(n1029) );
  MXI2X4 U1297 ( .A(n2072), .B(n1027), .S0(n1648), .Y(n1138) );
  NAND2X8 U1298 ( .A(n1034), .B(n1031), .Y(n1519) );
  NAND2X6 U1299 ( .A(n1035), .B(n1654), .Y(n1034) );
  NAND3X6 U1300 ( .A(n1038), .B(n1037), .C(n1036), .Y(n1035) );
  NAND3X8 U1301 ( .A(n1991), .B(n1471), .C(n1992), .Y(n1037) );
  NAND3X8 U1302 ( .A(n1402), .B(n1401), .C(n1400), .Y(n1038) );
  AOI21X4 U1303 ( .A0(n1995), .A1(n1994), .B0(n1040), .Y(n1039) );
  CLKINVX6 U1304 ( .A(n1996), .Y(n1040) );
  NAND2X4 U1305 ( .A(n1176), .B(n1989), .Y(n1042) );
  CLKINVX6 U1306 ( .A(CNT3[2]), .Y(n1044) );
  CLKBUFX8 U1307 ( .A(n2061), .Y(n1045) );
  NAND2BX4 U1308 ( .AN(n2061), .B(n2060), .Y(n2050) );
  MXI2X4 U1309 ( .A(n2145), .B(n1046), .S0(n1790), .Y(n2172) );
  MXI2X4 U1310 ( .A(n2145), .B(n1046), .S0(n1791), .Y(n2265) );
  CLKINVX6 U1311 ( .A(n1045), .Y(n1046) );
  MXI2X4 U1312 ( .A(n1048), .B(n1047), .S0(n1074), .Y(n2061) );
  CLKINVX6 U1313 ( .A(n1220), .Y(n1047) );
  CLKINVX6 U1314 ( .A(n669), .Y(n1048) );
  CLKINVX20 U1320 ( .A(n610), .Y(n1052) );
  NAND2X8 U1322 ( .A(n1411), .B(n1054), .Y(n1053) );
  INVX6 U1323 ( .A(n1055), .Y(n1054) );
  OR2X8 U1325 ( .A(n2594), .B(n611), .Y(n1056) );
  INVXL U1327 ( .A(n1931), .Y(n1974) );
  NOR2X8 U1328 ( .A(n1975), .B(n1931), .Y(n1513) );
  NAND2X8 U1329 ( .A(n1972), .B(n1932), .Y(n1515) );
  INVX12 U1330 ( .A(n1072), .Y(n1220) );
  NAND2X8 U1331 ( .A(n2043), .B(CNT5[4]), .Y(n1289) );
  NAND2X6 U1332 ( .A(n2248), .B(CNT6[3]), .Y(n2117) );
  INVX20 U1333 ( .A(n2123), .Y(n1082) );
  NAND2X4 U1334 ( .A(n2247), .B(CNT6[4]), .Y(n1631) );
  OR2X1 U1335 ( .A(n1323), .B(n1006), .Y(n1058) );
  OR2X4 U1336 ( .A(n2179), .B(n2084), .Y(n1059) );
  OR2X8 U1337 ( .A(n1663), .B(n1662), .Y(n1061) );
  INVX3 U1338 ( .A(n1590), .Y(n1063) );
  BUFX8 U1339 ( .A(n2000), .Y(n1064) );
  INVXL U1340 ( .A(n1233), .Y(n1929) );
  NOR2X4 U1341 ( .A(n2406), .B(n2407), .Y(n1543) );
  MXI2XL U1342 ( .A(n950), .B(n2089), .S0(n1330), .Y(n1777) );
  OR2X4 U1343 ( .A(n2171), .B(n2172), .Y(n1583) );
  MX2X8 U1344 ( .A(n950), .B(n2089), .S0(n1076), .Y(n2297) );
  CLKBUFX6 U1345 ( .A(n2091), .Y(n1219) );
  NAND2X8 U1346 ( .A(n1630), .B(n1425), .Y(n1424) );
  NAND2X6 U1347 ( .A(n1987), .B(n2088), .Y(n1986) );
  INVX6 U1348 ( .A(n2196), .Y(n1299) );
  MXI2X6 U1349 ( .A(n2614), .B(n2615), .S0(n1802), .Y(\com[4][6] ) );
  NAND3X8 U1351 ( .A(n2236), .B(n2235), .C(n2421), .Y(n2237) );
  MXI2X8 U1352 ( .A(n2597), .B(n1410), .S0(n1802), .Y(\com[4][2] ) );
  MXI2X8 U1355 ( .A(n2435), .B(n1444), .S0(n1802), .Y(\com[4][4] ) );
  MXI2X2 U1356 ( .A(n2624), .B(n2623), .S0(n1352), .Y(n1457) );
  AND2X6 U1357 ( .A(n1612), .B(n1616), .Y(n1090) );
  CLKINVX3 U1361 ( .A(n1525), .Y(n1087) );
  NAND2X4 U1362 ( .A(n2046), .B(n1970), .Y(n1269) );
  INVX1 U1363 ( .A(n2069), .Y(n2082) );
  CLKINVX2 U1364 ( .A(n1976), .Y(n1493) );
  NOR2X6 U1365 ( .A(n1602), .B(n1623), .Y(n1601) );
  INVX4 U1366 ( .A(n1779), .Y(n2239) );
  NAND2X8 U1367 ( .A(n2217), .B(n2387), .Y(n2218) );
  INVX6 U1368 ( .A(n1319), .Y(n2214) );
  INVX1 U1369 ( .A(n975), .Y(n2279) );
  NAND2X6 U1370 ( .A(n1762), .B(n1138), .Y(n1584) );
  MXI2X4 U1371 ( .A(n2298), .B(n1777), .S0(n1331), .Y(\com[2][2] ) );
  CLKMX2X6 U1372 ( .A(n2045), .B(n668), .S0(n1625), .Y(n1073) );
  AND2XL U1373 ( .A(n1006), .B(n2533), .Y(n2537) );
  NAND2X8 U1374 ( .A(n1220), .B(CNT5[2]), .Y(n2010) );
  MXI2X6 U1375 ( .A(n1329), .B(CNT5[5]), .S0(n1625), .Y(n1764) );
  CLKINVX1 U1376 ( .A(n1620), .Y(n1067) );
  CLKAND2X2 U1377 ( .A(n2614), .B(n2419), .Y(n1102) );
  NAND2X6 U1378 ( .A(n1930), .B(n657), .Y(n1903) );
  INVX6 U1379 ( .A(n1930), .Y(n1916) );
  INVX4 U1380 ( .A(n2248), .Y(n2120) );
  NAND3X6 U1381 ( .A(n2126), .B(n1393), .C(n1392), .Y(n1560) );
  NAND3X6 U1382 ( .A(n2125), .B(n2124), .C(n1082), .Y(n1392) );
  NAND2X6 U1383 ( .A(n1595), .B(n1594), .Y(n1657) );
  INVX8 U1384 ( .A(n1792), .Y(n1793) );
  CLKAND2X12 U1385 ( .A(n2156), .B(n1060), .Y(n1775) );
  INVX16 U1386 ( .A(n1652), .Y(n1389) );
  INVX20 U1387 ( .A(n1659), .Y(n1792) );
  BUFX16 U1388 ( .A(n1691), .Y(n1267) );
  MXI2X6 U1389 ( .A(n2090), .B(n1219), .S0(n1499), .Y(n2171) );
  NAND2X8 U1390 ( .A(n1558), .B(n1110), .Y(n1300) );
  CLKAND2X12 U1391 ( .A(n2156), .B(n1776), .Y(n2153) );
  INVX3 U1392 ( .A(n1801), .Y(n1146) );
  INVX4 U1393 ( .A(n1566), .Y(n2103) );
  INVX8 U1394 ( .A(n2084), .Y(n2180) );
  NAND2X4 U1395 ( .A(n1661), .B(n1660), .Y(n1426) );
  NOR2X8 U1396 ( .A(n2102), .B(n2398), .Y(n1277) );
  NOR2X8 U1397 ( .A(n1068), .B(n1273), .Y(n1545) );
  AND2X8 U1398 ( .A(n1773), .B(n2213), .Y(n1538) );
  INVX6 U1399 ( .A(n1338), .Y(n2136) );
  NAND2X6 U1400 ( .A(n2136), .B(n682), .Y(n2122) );
  NAND3X6 U1401 ( .A(n1530), .B(n2126), .C(n1532), .Y(n1562) );
  INVX6 U1402 ( .A(n2059), .Y(n2135) );
  NAND2X6 U1403 ( .A(n1477), .B(n1478), .Y(n2063) );
  AND2X6 U1404 ( .A(n2210), .B(n2411), .Y(n1069) );
  OR2X8 U1405 ( .A(n1625), .B(n669), .Y(n1679) );
  MXI2X8 U1406 ( .A(CNT5[4]), .B(n2113), .S0(n1789), .Y(n2139) );
  INVX20 U1407 ( .A(n1624), .Y(n1625) );
  AOI211X2 U1408 ( .A0(n2366), .A1(\com[2][1] ), .B0(n2355), .C0(n2354), .Y(
        n2360) );
  NAND2X8 U1409 ( .A(n1559), .B(n1104), .Y(n1178) );
  NOR2X6 U1410 ( .A(n1544), .B(n1543), .Y(n1534) );
  NOR2X6 U1411 ( .A(n2389), .B(n2390), .Y(n1537) );
  MXI2XL U1412 ( .A(n2535), .B(n1067), .S0(n2534), .Y(n2541) );
  NOR3X6 U1413 ( .A(n1757), .B(n1691), .C(n1565), .Y(n1564) );
  NOR2X6 U1414 ( .A(n1757), .B(n1691), .Y(n1286) );
  BUFX20 U1415 ( .A(n2661), .Y(n1803) );
  INVXL U1416 ( .A(n2210), .Y(n2412) );
  NOR2X6 U1417 ( .A(n2210), .B(n2411), .Y(n1544) );
  INVX6 U1418 ( .A(n2230), .Y(n2410) );
  CLKBUFX2 U1419 ( .A(n2217), .Y(n1142) );
  INVX12 U1420 ( .A(n2414), .Y(n2229) );
  INVXL U1421 ( .A(n2229), .Y(n1071) );
  NAND2X6 U1422 ( .A(n1978), .B(n1934), .Y(n1512) );
  AND2X4 U1423 ( .A(n2069), .B(n2081), .Y(n1404) );
  NAND2X8 U1424 ( .A(n1406), .B(n1404), .Y(n1400) );
  MX2X8 U1425 ( .A(n2009), .B(CNT4[2]), .S0(n1786), .Y(n1072) );
  INVX20 U1426 ( .A(n1421), .Y(n1638) );
  INVX12 U1427 ( .A(n1762), .Y(n1629) );
  CLKBUFX6 U1428 ( .A(n1662), .Y(n1563) );
  MXI2X4 U1429 ( .A(n2244), .B(n2402), .S0(n979), .Y(\com[3][7] ) );
  INVX3 U1430 ( .A(n1609), .Y(n1928) );
  NAND2X4 U1431 ( .A(n1379), .B(n1290), .Y(n2064) );
  INVX12 U1432 ( .A(n1195), .Y(n1648) );
  NAND3X6 U1433 ( .A(n1497), .B(n1495), .C(n1496), .Y(n1075) );
  BUFX12 U1434 ( .A(n1074), .Y(n1323) );
  INVX16 U1435 ( .A(n1792), .Y(n1076) );
  NAND2X8 U1436 ( .A(n2413), .B(n2229), .Y(n2231) );
  NAND2X4 U1437 ( .A(n1923), .B(n663), .Y(n1900) );
  BUFX16 U1438 ( .A(n1343), .Y(n1325) );
  NOR2X6 U1439 ( .A(n1194), .B(n1167), .Y(n1377) );
  NAND2X6 U1440 ( .A(n2059), .B(n1764), .Y(n2062) );
  MXI2X6 U1441 ( .A(CNT4[7]), .B(n1318), .S0(n1356), .Y(n2038) );
  CLKBUFX4 U1442 ( .A(n1071), .Y(n1296) );
  CLKAND2X12 U1443 ( .A(n1756), .B(n1319), .Y(n2198) );
  OAI2BB1X4 U1444 ( .A0N(n1221), .A1N(n1625), .B0(n1679), .Y(n2118) );
  OR2X4 U1445 ( .A(n1003), .B(n1760), .Y(n1248) );
  INVX8 U1446 ( .A(n1968), .Y(n1525) );
  NAND2X8 U1447 ( .A(n1606), .B(n1617), .Y(n1938) );
  NAND2X6 U1448 ( .A(n1065), .B(n1977), .Y(n1606) );
  NAND2X4 U1449 ( .A(n2292), .B(n2293), .Y(n2177) );
  CLKINVX4 U1450 ( .A(n2071), .Y(n1077) );
  INVX6 U1451 ( .A(n1077), .Y(n1078) );
  INVX4 U1452 ( .A(n2198), .Y(n2199) );
  NAND2X8 U1453 ( .A(n1224), .B(n1009), .Y(n1690) );
  INVX6 U1454 ( .A(n2139), .Y(n2071) );
  AND2X8 U1455 ( .A(n2139), .B(n2070), .Y(n1419) );
  NOR2X6 U1456 ( .A(n2297), .B(n2298), .Y(n2175) );
  MXI2X4 U1457 ( .A(n2116), .B(n665), .S0(n1789), .Y(n2141) );
  NAND2X4 U1458 ( .A(n2052), .B(n1954), .Y(n1311) );
  INVX8 U1459 ( .A(n1771), .Y(n2072) );
  NOR2X8 U1460 ( .A(n1428), .B(n1551), .Y(n1550) );
  MXI2X4 U1461 ( .A(n671), .B(n2115), .S0(n1323), .Y(n2150) );
  NAND2X8 U1462 ( .A(n1437), .B(n1436), .Y(n1785) );
  NAND2X8 U1463 ( .A(n1437), .B(n1436), .Y(n1137) );
  MXI2X4 U1464 ( .A(n2273), .B(n1291), .S0(n979), .Y(\com[3][6] ) );
  NAND2X6 U1465 ( .A(n1773), .B(n2213), .Y(n1272) );
  CLKBUFX2 U1466 ( .A(n1773), .Y(n1293) );
  INVX12 U1467 ( .A(n2233), .Y(n2413) );
  NAND2X6 U1468 ( .A(n2160), .B(n2159), .Y(n1571) );
  NOR2X6 U1469 ( .A(n2275), .B(n2405), .Y(n2205) );
  CLKINVX1 U1470 ( .A(n2419), .Y(n2273) );
  MX2X6 U1471 ( .A(n1080), .B(n2118), .S0(n1569), .Y(n2174) );
  CLKINVX20 U1472 ( .A(n685), .Y(n1080) );
  INVX8 U1473 ( .A(n2102), .Y(n1321) );
  MXI2X6 U1474 ( .A(n1301), .B(n2189), .S0(n1792), .Y(n1757) );
  NAND2X8 U1475 ( .A(n1552), .B(n1632), .Y(n1497) );
  MXI2X4 U1476 ( .A(n1527), .B(n1988), .S0(n1582), .Y(n1081) );
  MXI2X6 U1477 ( .A(n1774), .B(n2086), .S0(n1582), .Y(n2084) );
  NAND2X8 U1478 ( .A(n2147), .B(n2258), .Y(n1578) );
  INVX6 U1479 ( .A(n1760), .Y(n1408) );
  NOR2X4 U1480 ( .A(n2092), .B(n1760), .Y(n1428) );
  INVX3 U1481 ( .A(n1094), .Y(n1083) );
  NAND2X6 U1482 ( .A(n2392), .B(n1521), .Y(n1139) );
  AOI21X4 U1483 ( .A0(n1082), .A1(n1083), .B0(n1531), .Y(n1530) );
  NAND2X6 U1484 ( .A(n2236), .B(n2235), .Y(n2228) );
  MXI2X6 U1485 ( .A(n2226), .B(n1759), .S0(n1639), .Y(n2419) );
  NAND3X8 U1486 ( .A(n2065), .B(n1418), .C(n2063), .Y(n1378) );
  INVXL U1487 ( .A(n2134), .Y(n1084) );
  INVX3 U1488 ( .A(n1084), .Y(n1085) );
  MXI2X8 U1489 ( .A(n1088), .B(n2044), .S0(n1673), .Y(n2070) );
  INVX6 U1490 ( .A(n1087), .Y(n1088) );
  CLKINVX1 U1491 ( .A(n1330), .Y(n1086) );
  NAND2X6 U1492 ( .A(n1072), .B(n669), .Y(n2017) );
  INVX4 U1493 ( .A(n2045), .Y(n2112) );
  NAND2X8 U1494 ( .A(n1787), .B(n1655), .Y(n1354) );
  BUFX20 U1495 ( .A(n1519), .Y(n1499) );
  NAND2X6 U1496 ( .A(n2056), .B(n665), .Y(n2021) );
  NAND3X8 U1497 ( .A(n2030), .B(n2028), .C(n2029), .Y(n2035) );
  NAND2X6 U1498 ( .A(n1433), .B(n1432), .Y(n1604) );
  NAND3X6 U1499 ( .A(n1958), .B(n1957), .C(n1951), .Y(n1688) );
  NAND2X2 U1500 ( .A(n1973), .B(n1758), .Y(n1958) );
  NAND2X6 U1501 ( .A(n2140), .B(n2071), .Y(n1480) );
  INVX12 U1502 ( .A(n1232), .Y(n2045) );
  OR2X4 U1503 ( .A(n2049), .B(n1976), .Y(n1956) );
  INVX20 U1504 ( .A(n1353), .Y(n1787) );
  NAND2X8 U1505 ( .A(n1548), .B(n1278), .Y(n1496) );
  INVX20 U1506 ( .A(n1242), .Y(n1324) );
  NAND2X6 U1507 ( .A(n2419), .B(n2418), .Y(n2235) );
  CLKBUFX6 U1508 ( .A(n2389), .Y(n1292) );
  BUFX8 U1509 ( .A(n2224), .Y(n1420) );
  MXI2X8 U1510 ( .A(n1168), .B(n2093), .S0(n1582), .Y(n2092) );
  MXI2X4 U1511 ( .A(CNT4[4]), .B(n2003), .S0(n1356), .Y(n1215) );
  NAND2X8 U1512 ( .A(n1949), .B(n673), .Y(n1918) );
  OR2X8 U1513 ( .A(n1609), .B(CNT3[5]), .Y(n1904) );
  NAND2X6 U1514 ( .A(n1904), .B(n1903), .Y(n1901) );
  AND2XL U1515 ( .A(n972), .B(n2513), .Y(n2518) );
  NAND2X6 U1516 ( .A(n1235), .B(n1324), .Y(n1884) );
  NAND2X4 U1517 ( .A(n1175), .B(n2062), .Y(n1370) );
  NAND4X8 U1518 ( .A(n1939), .B(n1070), .C(n1938), .D(n1515), .Y(n1596) );
  BUFX12 U1519 ( .A(n2088), .Y(n1288) );
  NAND2X8 U1521 ( .A(n2183), .B(n2092), .Y(n1626) );
  BUFX20 U1522 ( .A(n2183), .Y(n1760) );
  NAND2X6 U1523 ( .A(n1151), .B(CNT3[2]), .Y(n1150) );
  NAND2X8 U1524 ( .A(n1609), .B(CNT3[5]), .Y(n1506) );
  MXI2X8 U1525 ( .A(n2135), .B(n1216), .S0(n1790), .Y(n2183) );
  INVX1 U1526 ( .A(n1342), .Y(n1899) );
  MXI2X8 U1527 ( .A(n1925), .B(n1926), .S0(n1024), .Y(n1917) );
  MXI2X6 U1528 ( .A(n2003), .B(CNT4[4]), .S0(n1786), .Y(n2043) );
  MXI2X6 U1529 ( .A(n1013), .B(n1078), .S0(n1790), .Y(n2179) );
  MXI2X4 U1530 ( .A(CNT5[6]), .B(n2056), .S0(n1789), .Y(n2142) );
  INVX20 U1531 ( .A(n1625), .Y(n1789) );
  OR2X2 U1532 ( .A(n2402), .B(n2431), .Y(n1307) );
  INVXL U1533 ( .A(\com[2][6] ), .Y(n1450) );
  MXI2X4 U1534 ( .A(n656), .B(n1921), .S0(n1326), .Y(n1943) );
  INVX1 U1535 ( .A(n1950), .Y(n1983) );
  INVX4 U1536 ( .A(n2426), .Y(n1667) );
  NOR2X6 U1537 ( .A(n2043), .B(CNT5[4]), .Y(n2024) );
  INVX3 U1538 ( .A(n2034), .Y(n2109) );
  MXI2X4 U1539 ( .A(n1948), .B(n1092), .S0(n1339), .Y(n2081) );
  NAND2X6 U1540 ( .A(n2424), .B(n1665), .Y(n1165) );
  INVX3 U1541 ( .A(n1414), .Y(n2424) );
  MXI2X4 U1542 ( .A(n1653), .B(n2136), .S0(n1569), .Y(n2257) );
  CLKINVX1 U1543 ( .A(n682), .Y(n1653) );
  CLKAND2X8 U1544 ( .A(n1631), .B(n1108), .Y(n1093) );
  NOR2X4 U1545 ( .A(n2123), .B(n1094), .Y(n1394) );
  INVXL U1546 ( .A(n2213), .Y(n2384) );
  INVX1 U1547 ( .A(n2601), .Y(n2602) );
  INVX3 U1548 ( .A(n1410), .Y(n1412) );
  INVX3 U1549 ( .A(n1759), .Y(n2400) );
  NAND2X2 U1550 ( .A(n2307), .B(n2482), .Y(n2309) );
  INVX3 U1551 ( .A(n1308), .Y(n1444) );
  MXI2X4 U1552 ( .A(n2611), .B(n989), .S0(n1803), .Y(\com[4][5] ) );
  NOR2X1 U1553 ( .A(gray_data[2]), .B(n2915), .Y(n2917) );
  INVX12 U1554 ( .A(n1244), .Y(n1768) );
  MXI2X1 U1555 ( .A(n2249), .B(n686), .S0(n1797), .Y(\com[0][1] ) );
  INVXL U1556 ( .A(n1757), .Y(n2286) );
  MXI2X2 U1557 ( .A(n2256), .B(n1312), .S0(n1798), .Y(\com[1][6] ) );
  CLKINVX1 U1558 ( .A(\com[1][6] ), .Y(n2770) );
  MXI2X1 U1559 ( .A(n2246), .B(n681), .S0(n1797), .Y(\com[0][6] ) );
  CLKINVX1 U1560 ( .A(\com[0][7] ), .Y(n1346) );
  MXI2X1 U1561 ( .A(n2253), .B(n2252), .S0(n1798), .Y(\com[1][7] ) );
  NOR3BXL U1562 ( .AN(gray_data[2]), .B(gray_data[1]), .C(n2915), .Y(n2916) );
  NOR3X4 U1563 ( .A(n2915), .B(n1866), .C(n1865), .Y(n1875) );
  CLKINVX1 U1564 ( .A(gray_data[2]), .Y(n1866) );
  CLKAND2X3 U1565 ( .A(gray_data[0]), .B(n2916), .Y(n1864) );
  INVX1 U1566 ( .A(n2268), .Y(n2269) );
  MXI2X1 U1567 ( .A(n2250), .B(n687), .S0(n1797), .Y(\com[0][0] ) );
  INVX4 U1568 ( .A(CNT1[0]), .Y(n1203) );
  NOR2X4 U1569 ( .A(n1846), .B(gray_data[1]), .Y(n1836) );
  NOR2X4 U1570 ( .A(n1846), .B(n1865), .Y(n1855) );
  NOR2X6 U1571 ( .A(n1342), .B(n1241), .Y(n1883) );
  NOR2X4 U1572 ( .A(n1768), .B(n1236), .Y(n1876) );
  NAND2X6 U1573 ( .A(n1774), .B(n1985), .Y(n1405) );
  NAND2X4 U1574 ( .A(n2389), .B(n2390), .Y(n1539) );
  MXI2X2 U1575 ( .A(n2042), .B(n2041), .S0(n1673), .Y(n2054) );
  NAND2XL U1576 ( .A(n1946), .B(n1945), .Y(n1996) );
  INVXL U1577 ( .A(n1944), .Y(n1945) );
  MXI2X4 U1578 ( .A(n1092), .B(n1948), .S0(n1217), .Y(n2052) );
  NOR2X6 U1579 ( .A(n1282), .B(n1281), .Y(n1427) );
  INVX2 U1580 ( .A(n1662), .Y(n1660) );
  CLKINVX1 U1581 ( .A(n1996), .Y(n1998) );
  INVX3 U1582 ( .A(n1650), .Y(n1574) );
  INVX3 U1583 ( .A(n1312), .Y(n1573) );
  INVX2 U1584 ( .A(n2097), .Y(n1527) );
  NAND2XL U1585 ( .A(n1620), .B(n1325), .Y(n2528) );
  OR2XL U1586 ( .A(n1620), .B(n1325), .Y(n2529) );
  NOR2X4 U1587 ( .A(n1949), .B(n1618), .Y(n1591) );
  NAND2XL U1588 ( .A(n1997), .B(n1998), .Y(n2106) );
  INVX3 U1589 ( .A(n2060), .Y(n2145) );
  INVX2 U1590 ( .A(n2080), .Y(n1581) );
  INVX3 U1591 ( .A(n2168), .Y(n1222) );
  NAND2X1 U1592 ( .A(n2398), .B(n2397), .Y(n2431) );
  INVX3 U1593 ( .A(n2298), .Y(n2204) );
  INVX4 U1594 ( .A(n2031), .Y(n2032) );
  NAND2XL U1595 ( .A(n1323), .B(n2513), .Y(n2519) );
  NOR2XL U1596 ( .A(n974), .B(n1336), .Y(n2514) );
  MXI2XL U1597 ( .A(n2701), .B(n2494), .S0(n974), .Y(n2495) );
  BUFX16 U1598 ( .A(n2225), .Y(n1759) );
  MXI2X4 U1599 ( .A(n1757), .B(n2227), .S0(n1799), .Y(n2418) );
  CLKINVX1 U1600 ( .A(n2106), .Y(n2397) );
  INVXL U1601 ( .A(n2203), .Y(n2394) );
  INVX1 U1602 ( .A(n2291), .Y(n1520) );
  CLKINVX1 U1603 ( .A(n2431), .Y(n2619) );
  INVXL U1604 ( .A(n1314), .Y(n2408) );
  NAND3X6 U1605 ( .A(n1160), .B(n1159), .C(n1165), .Y(n1158) );
  MXI2XL U1606 ( .A(n2647), .B(n2551), .S0(n1780), .Y(n2558) );
  OR2X1 U1607 ( .A(n1620), .B(n2493), .Y(n2535) );
  MXI2XL U1608 ( .A(n2498), .B(n2497), .S0(n981), .Y(n2501) );
  INVXL U1609 ( .A(n1292), .Y(n2391) );
  MXI2X4 U1610 ( .A(n2394), .B(n1285), .S0(n1639), .Y(n2392) );
  CLKINVX2 U1611 ( .A(n1445), .Y(n1446) );
  NAND4BX1 U1612 ( .AN(gray_data[3]), .B(gray_valid), .C(n2918), .D(n2919), 
        .Y(n2915) );
  MXI2X1 U1613 ( .A(n1686), .B(n682), .S0(n1797), .Y(\com[0][5] ) );
  MXI2X1 U1614 ( .A(n2248), .B(n684), .S0(n1797), .Y(\com[0][3] ) );
  OAI22XL U1615 ( .A0(n2344), .A1(n2343), .B0(n804), .B1(n634), .Y(n2345) );
  NAND2X1 U1616 ( .A(gray_data[0]), .B(n2917), .Y(n1846) );
  CLKINVX1 U1617 ( .A(gray_data[1]), .Y(n1865) );
  INVX3 U1618 ( .A(n2311), .Y(n1664) );
  NAND2X1 U1619 ( .A(n2633), .B(n2862), .Y(n1482) );
  INVX8 U1620 ( .A(n1213), .Y(n1214) );
  CLKBUFX3 U1621 ( .A(n1845), .Y(n1783) );
  NOR3BXL U1622 ( .AN(n2917), .B(n1865), .C(gray_data[0]), .Y(n1845) );
  OR2X1 U1624 ( .A(n2951), .B(tree_mem_back[2]), .Y(n2929) );
  OAI2BB1X1 U1625 ( .A0N(n2350), .A1N(n1726), .B0(n2644), .Y(n2936) );
  AOI21X1 U1626 ( .A0(\com[2][6] ), .A1(n1449), .B0(n2364), .Y(n1448) );
  OAI22XL U1627 ( .A0(n2347), .A1(n2346), .B0(n802), .B1(n636), .Y(n2348) );
  NOR2X2 U1628 ( .A(n2929), .B(n1818), .Y(n2913) );
  NAND2X2 U1629 ( .A(n2644), .B(n2942), .Y(n2939) );
  NAND2BX1 U1630 ( .AN(\com[1][7] ), .B(\com[0][7] ), .Y(n1344) );
  AOI2BB2X1 U1631 ( .B0(\com[1][7] ), .B1(n1346), .A0N(n2770), .A1N(
        \com[0][6] ), .Y(n1345) );
  INVXL U1632 ( .A(n1323), .Y(n2668) );
  NAND2X1 U1633 ( .A(state[1]), .B(n1711), .Y(n3046) );
  CLKINVX1 U1634 ( .A(n2939), .Y(n2910) );
  NOR2X2 U1635 ( .A(n2951), .B(n1728), .Y(n2911) );
  NOR2X1 U1636 ( .A(n2322), .B(n1738), .Y(n2585) );
  CLKBUFX3 U1637 ( .A(n2330), .Y(n1781) );
  NAND2X2 U1638 ( .A(n2271), .B(n2912), .Y(n2282) );
  OR2X1 U1639 ( .A(n2929), .B(n1817), .Y(n2932) );
  NAND2BX1 U1640 ( .AN(n2927), .B(n1740), .Y(n2322) );
  NAND2BX1 U1642 ( .AN(n3046), .B(n1712), .Y(n2927) );
  CLKBUFX3 U1643 ( .A(n1827), .Y(n1782) );
  CLKBUFX2 U1644 ( .A(n1898), .Y(CNT1[3]) );
  CLKBUFX2 U1645 ( .A(n1198), .Y(CNT1[7]) );
  OAI21XL U1646 ( .A0(n1855), .A1(n663), .B0(n1853), .Y(n849) );
  OAI21XL U1647 ( .A0(n1836), .A1(n1205), .B0(n1830), .Y(n829) );
  OAI21XL U1648 ( .A0(n1836), .A1(n1766), .B0(n1829), .Y(n828) );
  OAI21XL U1649 ( .A0(n1836), .A1(n1230), .B0(n1835), .Y(n826) );
  OAI21XL U1650 ( .A0(n1836), .A1(n1324), .B0(n1831), .Y(n830) );
  OAI21XL U1651 ( .A0(n1836), .A1(n1171), .B0(n1828), .Y(n827) );
  CLKINVX1 U1652 ( .A(n1781), .Y(n1135) );
  OAI2BB1X1 U1653 ( .A0N(n2284), .A1N(N1141), .B0(n2277), .Y(n812) );
  OAI21XL U1654 ( .A0(n1875), .A1(n686), .B0(n1872), .Y(n872) );
  OAI21XL U1655 ( .A0(n1875), .A1(n685), .B0(n1871), .Y(n871) );
  OAI21XL U1656 ( .A0(n1875), .A1(n684), .B0(n1870), .Y(n870) );
  OAI21XL U1657 ( .A0(n1875), .A1(n682), .B0(n1868), .Y(n868) );
  OAI21XL U1658 ( .A0(n1864), .A1(n669), .B0(n1860), .Y(n855) );
  OAI21XL U1659 ( .A0(n1864), .A1(n668), .B0(n1859), .Y(n854) );
  OAI21XL U1660 ( .A0(n1864), .A1(n667), .B0(n1858), .Y(n853) );
  OAI21XL U1661 ( .A0(n1864), .A1(n666), .B0(n1857), .Y(n852) );
  OAI2BB1X1 U1662 ( .A0N(n2284), .A1N(N1140), .B0(n2278), .Y(n811) );
  OAI21XL U1663 ( .A0(n1836), .A1(n1203), .B0(n1834), .Y(n833) );
  OAI21XL U1664 ( .A0(n1855), .A1(n656), .B0(n1854), .Y(n842) );
  OAI21XL U1665 ( .A0(n1855), .A1(n657), .B0(n1847), .Y(n843) );
  OAI21XL U1666 ( .A0(n1855), .A1(n658), .B0(n1848), .Y(n844) );
  OAI21XL U1667 ( .A0(n1855), .A1(n659), .B0(n1849), .Y(n845) );
  OAI21XL U1668 ( .A0(n1855), .A1(n660), .B0(n1850), .Y(n846) );
  OAI21XL U1669 ( .A0(n1855), .A1(n661), .B0(n1851), .Y(n847) );
  OAI21XL U1670 ( .A0(n1855), .A1(n662), .B0(n1852), .Y(n848) );
  INVX4 U1671 ( .A(n2214), .Y(n1140) );
  INVX12 U1673 ( .A(n1756), .Y(n2287) );
  MXI2X4 U1674 ( .A(n1475), .B(n1476), .S0(n1325), .Y(n1092) );
  MXI2X4 U1675 ( .A(n664), .B(n2109), .S0(n1789), .Y(n2066) );
  INVX1 U1676 ( .A(n976), .Y(n2457) );
  BUFX3 U1677 ( .A(n2037), .Y(n1280) );
  INVXL U1678 ( .A(n2114), .Y(n2249) );
  INVX8 U1679 ( .A(n1391), .Y(n2247) );
  CLKINVX8 U1680 ( .A(n1476), .Y(CNT1[1]) );
  CLKINVX8 U1681 ( .A(n1475), .Y(CNT2[1]) );
  CLKBUFX2 U1682 ( .A(n1339), .Y(n1620) );
  CLKINVX12 U1683 ( .A(n1335), .Y(n1353) );
  INVX3 U1684 ( .A(n1521), .Y(n2393) );
  INVX3 U1685 ( .A(n954), .Y(n2256) );
  BUFX12 U1686 ( .A(n1799), .Y(n1331) );
  INVX4 U1687 ( .A(n1985), .Y(n2086) );
  INVX1 U1688 ( .A(n1798), .Y(n1265) );
  CLKBUFX8 U1689 ( .A(n1383), .Y(n1798) );
  INVX8 U1690 ( .A(n1207), .Y(n1208) );
  INVX12 U1691 ( .A(n1212), .Y(n1885) );
  INVX12 U1692 ( .A(n1885), .Y(CNT2[2]) );
  INVX12 U1693 ( .A(n1243), .Y(n1342) );
  INVX3 U1694 ( .A(n1899), .Y(n1476) );
  INVX6 U1695 ( .A(n2600), .Y(n2417) );
  BUFX12 U1696 ( .A(n1582), .Y(n1526) );
  INVX3 U1697 ( .A(\com[3][7] ), .Y(n2378) );
  OR2X8 U1698 ( .A(n2247), .B(CNT6[4]), .Y(n1094) );
  MXI2X4 U1699 ( .A(n661), .B(n1929), .S0(n1025), .Y(n1978) );
  CLKBUFX3 U1700 ( .A(n1063), .Y(n1318) );
  INVX3 U1701 ( .A(n1999), .Y(n1590) );
  INVX6 U1702 ( .A(n2201), .Y(n1565) );
  CLKINVX4 U1703 ( .A(n1241), .Y(n1475) );
  INVX1 U1704 ( .A(n2075), .Y(n2108) );
  INVX3 U1705 ( .A(\com[4][4] ), .Y(n2467) );
  AND2X2 U1706 ( .A(n2913), .B(n1726), .Y(n1095) );
  BUFX12 U1707 ( .A(n1137), .Y(n1326) );
  CLKBUFX3 U1708 ( .A(n1356), .Y(n1336) );
  INVX3 U1709 ( .A(n1971), .Y(n1932) );
  INVX3 U1710 ( .A(n2407), .Y(n1567) );
  CLKAND2X12 U1711 ( .A(n2620), .B(n2431), .Y(n1098) );
  OA22X2 U1712 ( .A0(\com[3][6] ), .A1(n635), .B0(\com[3][5] ), .B1(n634), .Y(
        n1099) );
  INVX1 U1713 ( .A(n1379), .Y(n1216) );
  MXI2X8 U1714 ( .A(n2404), .B(n1284), .S0(n1313), .Y(n1100) );
  INVX4 U1715 ( .A(\com[3][6] ), .Y(n1449) );
  INVX4 U1716 ( .A(n1179), .Y(n1177) );
  INVX3 U1717 ( .A(n2181), .Y(n2260) );
  INVX8 U1718 ( .A(n1658), .Y(\com[2][5] ) );
  CLKMX2X4 U1719 ( .A(n2287), .B(n1140), .S0(n1331), .Y(n1658) );
  INVX3 U1720 ( .A(n2597), .Y(n1672) );
  MXI2X4 U1721 ( .A(n1293), .B(n2384), .S0(n1796), .Y(n2611) );
  BUFX12 U1722 ( .A(n1767), .Y(CNT1[5]) );
  INVX3 U1724 ( .A(n2131), .Y(n1481) );
  AND2X4 U1725 ( .A(n1270), .B(n1944), .Y(n1103) );
  INVX6 U1726 ( .A(n2435), .Y(n2612) );
  CLKAND2X12 U1727 ( .A(n2105), .B(n2106), .Y(n1104) );
  CLKINVX1 U1728 ( .A(n2399), .Y(n2226) );
  MXI2X2 U1729 ( .A(n2097), .B(n2096), .S0(n1788), .Y(n2399) );
  OA21X4 U1730 ( .A0(n1949), .A1(n673), .B0(n672), .Y(n1105) );
  INVX1 U1731 ( .A(n2066), .Y(n2132) );
  OR2X6 U1732 ( .A(n2159), .B(n2251), .Y(n2201) );
  CLKINVX1 U1733 ( .A(n2390), .Y(n1540) );
  MXI2X6 U1734 ( .A(n977), .B(n1296), .S0(n1313), .Y(\com[3][3] ) );
  AND2X2 U1735 ( .A(\com[3][6] ), .B(n1450), .Y(n1107) );
  OR2X4 U1736 ( .A(n2114), .B(n686), .Y(n1108) );
  AND3X8 U1737 ( .A(n1578), .B(n2148), .C(n1645), .Y(n1109) );
  CLKAND2X12 U1738 ( .A(n2103), .B(n2398), .Y(n1110) );
  NAND2X4 U1739 ( .A(n2430), .B(n2619), .Y(n2426) );
  INVX4 U1740 ( .A(n2090), .Y(n1492) );
  CLKINVX1 U1741 ( .A(n2077), .Y(n2107) );
  OR2X4 U1742 ( .A(n2066), .B(n2131), .Y(n2077) );
  INVXL U1743 ( .A(n1988), .Y(n2096) );
  INVXL U1744 ( .A(n2290), .Y(n1523) );
  INVX3 U1745 ( .A(n2055), .Y(n2133) );
  AND2X4 U1746 ( .A(n2234), .B(n2402), .Y(n1111) );
  MXI2X2 U1747 ( .A(n2285), .B(n1565), .S0(n1780), .Y(\com[2][7] ) );
  CLKINVX1 U1748 ( .A(\com[2][7] ), .Y(n2485) );
  INVX3 U1749 ( .A(n1770), .Y(CNT1[2]) );
  OR2X1 U1750 ( .A(n2938), .B(n614), .Y(n1112) );
  INVX8 U1751 ( .A(n1208), .Y(CNT2[5]) );
  INVX16 U1752 ( .A(n1526), .Y(n1788) );
  MX2XL U1753 ( .A(n2660), .B(n2659), .S0(n1352), .Y(n1117) );
  MX2XL U1754 ( .A(n2573), .B(n2574), .S0(n1012), .Y(n1119) );
  MXI2X1 U1755 ( .A(n2517), .B(n2516), .S0(n1796), .Y(n1120) );
  NOR2X2 U1756 ( .A(n2709), .B(n2729), .Y(n1134) );
  INVX12 U1757 ( .A(n1331), .Y(n1780) );
  OA22X4 U1760 ( .A0(n1100), .A1(n631), .B0(\com[3][3] ), .B1(n632), .Y(n2299)
         );
  INVX16 U1768 ( .A(n1467), .Y(\com[3][1] ) );
  NAND2X6 U1769 ( .A(n1186), .B(n1099), .Y(n2316) );
  NOR3X4 U1770 ( .A(n1801), .B(n1291), .C(n2623), .Y(n2403) );
  AOI2BB1X4 U1773 ( .A0N(n2360), .A1N(n2359), .B0(n2358), .Y(n2363) );
  MXI2X4 U1775 ( .A(n2328), .B(n3246), .S0(n3127), .Y(n808) );
  INVX8 U1776 ( .A(\com[3][3] ), .Y(n2371) );
  MXI2X4 U1778 ( .A(n2329), .B(n3245), .S0(n3127), .Y(n807) );
  CLKBUFX3 U1780 ( .A(\com[4][1] ), .Y(n1445) );
  INVX2 U1784 ( .A(\com[4][2] ), .Y(n2461) );
  OAI21X4 U1786 ( .A0(n1352), .A1(n2604), .B0(n793), .Y(n2605) );
  INVXL U1788 ( .A(\com[4][6] ), .Y(n2452) );
  BUFX4 U1790 ( .A(n1922), .Y(n1228) );
  NAND2X4 U1791 ( .A(n1342), .B(n1241), .Y(n1881) );
  CLKINVX16 U1792 ( .A(n1586), .Y(n1249) );
  NAND2X6 U1793 ( .A(n1233), .B(n661), .Y(n1505) );
  CLKBUFX6 U1794 ( .A(n1784), .Y(n1343) );
  NAND2X2 U1795 ( .A(n1609), .B(CNT3[5]), .Y(n1906) );
  BUFX12 U1796 ( .A(n1249), .Y(n1149) );
  MXI2X8 U1798 ( .A(n978), .B(n1283), .S0(n1313), .Y(\com[3][5] ) );
  NOR2X1 U1800 ( .A(n1100), .B(n2353), .Y(n2354) );
  AOI211X4 U1801 ( .A0(\com[3][1] ), .A1(n2352), .B0(n2351), .C0(\com[3][0] ), 
        .Y(n2355) );
  OAI22X1 U1805 ( .A0(n2371), .A1(\com[2][3] ), .B0(n2367), .B1(\com[2][2] ), 
        .Y(n2359) );
  INVX4 U1806 ( .A(\com[4][5] ), .Y(n2468) );
  INVX1 U1809 ( .A(n3139), .Y(n2466) );
  NAND2X8 U1811 ( .A(n1441), .B(n1440), .Y(n1436) );
  INVX8 U1812 ( .A(n2265), .Y(n2173) );
  MXI2X1 U1813 ( .A(n2265), .B(n2264), .S0(n1798), .Y(\com[1][2] ) );
  CLKINVX4 U1814 ( .A(n2082), .Y(n1579) );
  CLKBUFX2 U1815 ( .A(n1911), .Y(n1340) );
  AND2X4 U1816 ( .A(n1922), .B(CNT3[1]), .Y(n1507) );
  NAND2X8 U1817 ( .A(n1911), .B(CNT3[4]), .Y(n1509) );
  INVX8 U1818 ( .A(n2603), .Y(n2598) );
  INVX12 U1819 ( .A(n2222), .Y(n1772) );
  AOI21X4 U1820 ( .A0(n2206), .A1(n1139), .B0(n2205), .Y(n2221) );
  BUFX16 U1821 ( .A(n2215), .Y(n1756) );
  AND2X8 U1822 ( .A(n1310), .B(n1480), .Y(n2065) );
  NAND2X8 U1823 ( .A(n1669), .B(n1381), .Y(n1668) );
  OAI21X4 U1824 ( .A0(n2423), .A1(n1667), .B0(n1665), .Y(n1159) );
  MXI2X4 U1825 ( .A(n1304), .B(n2416), .S0(n1796), .Y(n2451) );
  MXI2X8 U1826 ( .A(n1140), .B(n2287), .S0(n1799), .Y(n2222) );
  NAND2X8 U1827 ( .A(n1755), .B(n2188), .Y(n2076) );
  NAND2X8 U1828 ( .A(n2320), .B(n2319), .Y(n1141) );
  CLKAND2X12 U1829 ( .A(n2432), .B(n1381), .Y(n1155) );
  CLKAND2X12 U1830 ( .A(n2428), .B(n1409), .Y(n1157) );
  NAND3X8 U1831 ( .A(n1157), .B(n1156), .C(n1155), .Y(n1148) );
  NOR2X8 U1832 ( .A(n1670), .B(n1098), .Y(n1416) );
  NAND2X4 U1833 ( .A(n2624), .B(n2614), .Y(n2429) );
  INVX4 U1834 ( .A(n2432), .Y(n1305) );
  INVX6 U1835 ( .A(n2451), .Y(n2595) );
  OR2X8 U1836 ( .A(n2613), .B(n2427), .Y(n1671) );
  NOR2X8 U1837 ( .A(n1143), .B(n1305), .Y(n1164) );
  NAND2X6 U1840 ( .A(n2425), .B(n1414), .Y(n2624) );
  NAND2X8 U1841 ( .A(n1146), .B(n1145), .Y(n1414) );
  INVX8 U1842 ( .A(n1291), .Y(n1145) );
  NOR2X8 U1843 ( .A(n2403), .B(n1306), .Y(n1409) );
  NAND2X4 U1844 ( .A(n1309), .B(n2396), .Y(n1163) );
  BUFX4 U1845 ( .A(n2450), .Y(n1147) );
  BUFX8 U1846 ( .A(n2445), .Y(n1410) );
  NAND4X8 U1847 ( .A(n1161), .B(n1148), .C(n1158), .D(n1154), .Y(n2661) );
  AND2X8 U1848 ( .A(n1508), .B(n1150), .Y(n1502) );
  MXI2X4 U1849 ( .A(CNT1[2]), .B(CNT2[2]), .S0(n1149), .Y(n1151) );
  NAND2X4 U1850 ( .A(n1902), .B(CNT3[3]), .Y(n1508) );
  MXI2X4 U1851 ( .A(n1898), .B(n1235), .S0(n1249), .Y(n1902) );
  NAND3BX4 U1852 ( .AN(n1671), .B(n2429), .C(n2428), .Y(n1154) );
  NAND2X8 U1853 ( .A(n1415), .B(n2433), .Y(n1156) );
  NAND2X6 U1854 ( .A(n1416), .B(n2420), .Y(n1160) );
  NAND3X8 U1855 ( .A(n1164), .B(n1163), .C(n1162), .Y(n1161) );
  NOR2X8 U1856 ( .A(n2598), .B(n2417), .Y(n1166) );
  NAND3X4 U1857 ( .A(n1175), .B(n2062), .C(n2066), .Y(n1167) );
  BUFX4 U1858 ( .A(n2094), .Y(n1168) );
  MXI2X4 U1859 ( .A(n1001), .B(n1974), .S0(n1339), .Y(n2093) );
  NOR2X8 U1860 ( .A(n1501), .B(n1169), .Y(n1435) );
  NAND3X8 U1861 ( .A(n1904), .B(n1903), .C(CNT3[7]), .Y(n1169) );
  CLKAND2X12 U1862 ( .A(n1506), .B(n1905), .Y(n1501) );
  NAND2X6 U1863 ( .A(n2260), .B(n2182), .Y(n1577) );
  NAND4X8 U1864 ( .A(n1170), .B(n1627), .C(n1584), .D(n1626), .Y(n1554) );
  NAND2X8 U1865 ( .A(n1275), .B(n1274), .Y(n1170) );
  BUFX8 U1866 ( .A(n1768), .Y(n1171) );
  CLKINVX16 U1867 ( .A(n1227), .Y(n1766) );
  INVXL U1868 ( .A(n1204), .Y(n1205) );
  NAND2BX4 U1869 ( .AN(n1204), .B(n1210), .Y(n1172) );
  MXI2X4 U1870 ( .A(n1398), .B(n957), .S0(n1367), .Y(n2088) );
  INVX8 U1871 ( .A(n1764), .Y(n1379) );
  INVX3 U1872 ( .A(n1229), .Y(n1174) );
  NOR2X6 U1873 ( .A(n1174), .B(n1238), .Y(n1878) );
  MXI2X4 U1874 ( .A(n1088), .B(n2044), .S0(n1360), .Y(n1473) );
  MXI2X4 U1875 ( .A(n1981), .B(n1982), .S0(n1360), .Y(n2097) );
  MXI2X4 U1876 ( .A(n980), .B(n2058), .S0(n1360), .Y(n2073) );
  NAND2X8 U1877 ( .A(n2142), .B(n2073), .Y(n1175) );
  NAND2X8 U1878 ( .A(n2097), .B(n1988), .Y(n1176) );
  MXI2X4 U1879 ( .A(n1002), .B(n1177), .S0(n1360), .Y(n1290) );
  INVX4 U1880 ( .A(n1001), .Y(n1655) );
  NAND3X6 U1881 ( .A(n1378), .B(n1380), .C(n1369), .Y(n1368) );
  AND2X8 U1882 ( .A(n2179), .B(n2084), .Y(n1553) );
  NAND2X8 U1883 ( .A(n1178), .B(n1300), .Y(n1421) );
  CLKBUFX4 U1884 ( .A(n2048), .Y(n1179) );
  INVX8 U1885 ( .A(n1893), .Y(n1334) );
  MXI2X4 U1886 ( .A(n2085), .B(n2084), .S0(n1494), .Y(n2210) );
  NOR2X6 U1887 ( .A(n1180), .B(n1544), .Y(n1533) );
  AND2X8 U1888 ( .A(n1763), .B(n2415), .Y(n1180) );
  MXI2X4 U1889 ( .A(n1014), .B(n1762), .S0(n1494), .Y(n1763) );
  NAND2X4 U1890 ( .A(n1181), .B(n2318), .Y(n2319) );
  NAND2X4 U1891 ( .A(n2316), .B(n1182), .Y(n1181) );
  NOR2BX4 U1892 ( .AN(n2304), .B(n1183), .Y(n1182) );
  NAND2X4 U1893 ( .A(n2317), .B(n1184), .Y(n1183) );
  NOR2X6 U1894 ( .A(\com[3][7] ), .B(n1185), .Y(n1184) );
  NAND2X4 U1895 ( .A(n2484), .B(n2485), .Y(n1185) );
  NAND2X1 U1896 ( .A(n1188), .B(n1189), .Y(\com[0][2] ) );
  CLKINVX1 U1897 ( .A(n1797), .Y(n1190) );
  NAND2X1 U1898 ( .A(n1797), .B(CNT6[2]), .Y(n1188) );
  NAND2X1 U1899 ( .A(n2118), .B(n1190), .Y(n1189) );
  CLKBUFX4 U1900 ( .A(n2842), .Y(n1797) );
  MX2XL U1901 ( .A(n2258), .B(n1015), .S0(n1798), .Y(\com[1][5] ) );
  INVXL U1902 ( .A(\com[1][5] ), .Y(n1191) );
  NOR2XL U1903 ( .A(n2756), .B(\com[0][2] ), .Y(n2759) );
  INVXL U1904 ( .A(\com[0][2] ), .Y(n2753) );
  NOR2XL U1905 ( .A(n1191), .B(n2750), .Y(n2761) );
  CLKINVX2 U1906 ( .A(n1171), .Y(CNT1[6]) );
  CLKINVX2 U1907 ( .A(n2223), .Y(n1192) );
  CLKINVX6 U1908 ( .A(n2409), .Y(n2223) );
  INVX6 U1909 ( .A(n1513), .Y(n1939) );
  OR2X8 U1910 ( .A(n1922), .B(CNT3[1]), .Y(n1231) );
  CLKBUFX6 U1911 ( .A(n1288), .Y(n1317) );
  NAND2X6 U1912 ( .A(n1387), .B(n1385), .Y(n1193) );
  NAND2X8 U1913 ( .A(n2137), .B(n2138), .Y(n1569) );
  NOR2X4 U1914 ( .A(n1079), .B(n1573), .Y(n1572) );
  NAND2X4 U1915 ( .A(n2138), .B(n2137), .Y(n2842) );
  INVX6 U1916 ( .A(n1555), .Y(n1637) );
  INVX4 U1917 ( .A(n2160), .Y(n2161) );
  NAND2X8 U1918 ( .A(n1982), .B(n2058), .Y(n1961) );
  INVX20 U1919 ( .A(n1347), .Y(n1586) );
  AND2X8 U1920 ( .A(n2196), .B(n2195), .Y(n1425) );
  INVX4 U1921 ( .A(n1284), .Y(n1413) );
  CLKBUFX6 U1922 ( .A(n2165), .Y(n1337) );
  OAI21XL U1923 ( .A0(n1836), .A1(n1476), .B0(n1833), .Y(n832) );
  INVX1 U1924 ( .A(n1239), .Y(n1196) );
  NOR3X6 U1925 ( .A(n1895), .B(n1894), .C(n1893), .Y(n1896) );
  NOR2X8 U1926 ( .A(n1235), .B(n1324), .Y(n1888) );
  NAND2X6 U1927 ( .A(n2035), .B(n1685), .Y(n1224) );
  INVX6 U1928 ( .A(n1235), .Y(n1199) );
  NOR2X6 U1929 ( .A(n647), .B(n1213), .Y(n1882) );
  NAND2X6 U1930 ( .A(n1334), .B(n1892), .Y(n1201) );
  CLKBUFX2 U1931 ( .A(n1229), .Y(n1198) );
  INVX3 U1932 ( .A(n1199), .Y(CNT2[3]) );
  INVX2 U1933 ( .A(n1878), .Y(n1202) );
  NAND2X6 U1934 ( .A(n1202), .B(n1201), .Y(n1588) );
  NAND2X6 U1935 ( .A(n1897), .B(n1896), .Y(n1348) );
  CLKINVX12 U1936 ( .A(n1206), .Y(n1770) );
  CLKBUFX2 U1937 ( .A(n1196), .Y(CNT2[7]) );
  NOR2X4 U1938 ( .A(n1208), .B(n1767), .Y(n1894) );
  MXI2XL U1939 ( .A(n1770), .B(n1885), .S0(n1343), .Y(n1913) );
  INVXL U1940 ( .A(n1210), .Y(n1211) );
  OAI21XL U1941 ( .A0(n1836), .A1(n1770), .B0(n1832), .Y(n831) );
  NOR2X8 U1942 ( .A(n1766), .B(n1207), .Y(n1877) );
  CLKBUFX2 U1943 ( .A(n1210), .Y(CNT2[4]) );
  NOR2X8 U1944 ( .A(n1501), .B(n1901), .Y(n1439) );
  NOR2X4 U1945 ( .A(n1208), .B(n1767), .Y(n1245) );
  CLKBUFX2 U1946 ( .A(n1213), .Y(CNT2[0]) );
  MXI2X4 U1947 ( .A(CNT3[1]), .B(n1615), .S0(n1025), .Y(n1947) );
  INVX3 U1948 ( .A(n1917), .Y(n2003) );
  INVX6 U1949 ( .A(n2266), .Y(n2163) );
  MX2X4 U1950 ( .A(n2042), .B(n2041), .S0(n974), .Y(n1218) );
  CLKAND2X12 U1951 ( .A(n1986), .B(n1524), .Y(n1992) );
  CLKINVX2 U1952 ( .A(n2172), .Y(n2089) );
  INVX6 U1953 ( .A(n1980), .Y(n2094) );
  INVX1 U1954 ( .A(n1220), .Y(n1221) );
  INVX1 U1955 ( .A(n1222), .Y(n1223) );
  MXI2XL U1956 ( .A(n2260), .B(n2259), .S0(n1798), .Y(\com[1][4] ) );
  CLKBUFX2 U1957 ( .A(n1076), .Y(n1330) );
  CLKBUFX4 U1958 ( .A(n1763), .Y(n1304) );
  CLKBUFX6 U1959 ( .A(n2111), .Y(n1329) );
  NAND2X8 U1960 ( .A(n1505), .B(n1510), .Y(n1907) );
  NAND2X8 U1961 ( .A(n1927), .B(n660), .Y(n1510) );
  INVX16 U1962 ( .A(n1970), .Y(n2047) );
  CLKINVX4 U1963 ( .A(n1268), .Y(n1225) );
  CLKBUFX2 U1964 ( .A(n2051), .Y(n1268) );
  INVX4 U1965 ( .A(n2051), .Y(n2110) );
  NOR2X6 U1966 ( .A(n2047), .B(n1398), .Y(n1246) );
  OR2X6 U1967 ( .A(n1915), .B(CNT4[5]), .Y(n1518) );
  INVX4 U1968 ( .A(n1340), .Y(n1925) );
  INVX4 U1969 ( .A(n973), .Y(n2001) );
  BUFX20 U1970 ( .A(n1271), .Y(n1226) );
  BUFX16 U1971 ( .A(n2025), .Y(n1271) );
  NAND2X8 U1972 ( .A(n1986), .B(n1524), .Y(n1403) );
  OR2X6 U1973 ( .A(n951), .B(CNT5[3]), .Y(n1678) );
  INVX12 U1974 ( .A(n2046), .Y(n1398) );
  NOR3X4 U1975 ( .A(n1878), .B(n1877), .C(n1876), .Y(n1879) );
  INVX20 U1976 ( .A(n1766), .Y(n1767) );
  NAND3X8 U1977 ( .A(n2030), .B(n2018), .C(n2019), .Y(n2020) );
  BUFX20 U1978 ( .A(n2661), .Y(n1802) );
  BUFX16 U1979 ( .A(n1786), .Y(n1279) );
  AND3X8 U1980 ( .A(n2101), .B(n2100), .C(n1321), .Y(n1640) );
  NAND3X8 U1981 ( .A(n1363), .B(n1359), .C(n1362), .Y(n1358) );
  NAND3X8 U1982 ( .A(n1960), .B(n1687), .C(n1955), .Y(n1362) );
  INVX6 U1983 ( .A(n2013), .Y(n2111) );
  NAND2X6 U1984 ( .A(n1589), .B(n1588), .Y(n1587) );
  NOR2X4 U1985 ( .A(n1911), .B(CNT3[4]), .Y(n1905) );
  CLKINVX12 U1986 ( .A(n1586), .Y(n1784) );
  MXI2X4 U1987 ( .A(CNT1[1]), .B(CNT2[1]), .S0(n1784), .Y(n1922) );
  INVXL U1988 ( .A(n1198), .Y(n1230) );
  INVX4 U1989 ( .A(n1500), .Y(n1910) );
  AND2X8 U1990 ( .A(n1070), .B(n1515), .Y(n1327) );
  NAND2X4 U1991 ( .A(n1231), .B(n1900), .Y(n1504) );
  NAND2X6 U1992 ( .A(n2013), .B(CNT5[5]), .Y(n2025) );
  NAND2X4 U1993 ( .A(n2021), .B(n2022), .Y(n2015) );
  NOR2X8 U1994 ( .A(n1403), .B(n1407), .Y(n1402) );
  MXI2X4 U1995 ( .A(n964), .B(n676), .S0(n1786), .Y(n1232) );
  INVX12 U1996 ( .A(n1952), .Y(n2002) );
  NOR2X8 U1997 ( .A(n1266), .B(n2039), .Y(n1964) );
  CLKBUFX4 U1998 ( .A(n2405), .Y(n1284) );
  MXI2X4 U1999 ( .A(n2204), .B(n2297), .S0(n982), .Y(n2405) );
  AOI22X2 U2000 ( .A0(n633), .A1(\com[3][4] ), .B0(\com[3][5] ), .B1(n634), 
        .Y(n2302) );
  MXI2X4 U2001 ( .A(n1770), .B(n1885), .S0(n1149), .Y(n1233) );
  CLKINVX1 U2002 ( .A(CNT2[6]), .Y(n1234) );
  CLKBUFX2 U2003 ( .A(n1236), .Y(CNT2[6]) );
  INVXL U2004 ( .A(n1236), .Y(n1237) );
  INVXL U2005 ( .A(n1238), .Y(n1239) );
  CLKBUFX2 U2006 ( .A(n1204), .Y(CNT1[4]) );
  NAND2X8 U2007 ( .A(n1287), .B(n1599), .Y(n1316) );
  BUFX16 U2008 ( .A(n2288), .Y(n1761) );
  AOI2BB1X4 U2009 ( .A0N(n1215), .A1N(n1968), .B0(n1246), .Y(n1364) );
  NAND2X6 U2010 ( .A(n1509), .B(n1506), .Y(n1333) );
  CLKINVX2 U2011 ( .A(n2006), .Y(n2007) );
  NAND2X6 U2012 ( .A(n2158), .B(n2157), .Y(n1390) );
  INVX8 U2013 ( .A(n2224), .Y(n2386) );
  MXI2X4 U2014 ( .A(n2411), .B(n2412), .S0(n1639), .Y(n2409) );
  INVX8 U2015 ( .A(n2216), .Y(n2387) );
  NAND2X8 U2016 ( .A(n1629), .B(n1016), .Y(n1275) );
  CLKINVX8 U2017 ( .A(n1142), .Y(n1247) );
  NAND2X6 U2018 ( .A(n1539), .B(n1541), .Y(n1535) );
  NAND3X8 U2019 ( .A(n1533), .B(n2098), .C(n2099), .Y(n1641) );
  MXI2X2 U2020 ( .A(n2090), .B(n1219), .S0(n1526), .Y(n2407) );
  NAND2BX4 U2021 ( .AN(n1242), .B(n1235), .Y(n1886) );
  INVX4 U2022 ( .A(n1228), .Y(n1615) );
  INVXL U2023 ( .A(n1119), .Y(n1250) );
  MXI2X1 U2024 ( .A(n2503), .B(n2502), .S0(n1796), .Y(n2569) );
  AOI2BB2X2 U2025 ( .B0(n1265), .B1(n2577), .A0N(n2664), .A1N(n2695), .Y(n2709) );
  NAND2BX1 U2026 ( .AN(n2946), .B(state[2]), .Y(N202) );
  MXI2X4 U2027 ( .A(n968), .B(n1966), .S0(n1339), .Y(n2068) );
  INVXL U2028 ( .A(n1117), .Y(n1251) );
  OAI21X4 U2029 ( .A0(n2999), .A1(n2908), .B0(n1754), .Y(N686) );
  OAI211X4 U2030 ( .A0(n2739), .A1(n2737), .B0(n2581), .C0(n2580), .Y(N714) );
  OAI31X4 U2031 ( .A0(n2789), .A1(n2788), .A2(n2787), .B0(n2786), .Y(N658) );
  NAND2BXL U2032 ( .AN(n3058), .B(n2932), .Y(n728) );
  OAI211XL U2033 ( .A0(n1718), .A1(n3021), .B0(n1751), .C0(n3022), .Y(N667) );
  OAI211XL U2034 ( .A0(n1718), .A1(n2846), .B0(n2845), .C0(n2844), .Y(N723) );
  OAI211XL U2035 ( .A0(n1718), .A1(n3002), .B0(n3003), .C0(n3004), .Y(N681) );
  OAI211XL U2036 ( .A0(n3031), .A1(n1718), .B0(n3032), .C0(n3033), .Y(N653) );
  AOI2BB2XL U2037 ( .B0(n2899), .B1(n3069), .A0N(n3009), .A1N(n1733), .Y(n3017) );
  AOI2BB2XL U2038 ( .B0(n2898), .B1(n3069), .A0N(n3025), .A1N(n1733), .Y(n3030) );
  AOI2BB2XL U2039 ( .B0(n2905), .B1(n3069), .A0N(n2961), .A1N(n1714), .Y(n2976) );
  AOI2BB2XL U2040 ( .B0(n2905), .B1(n3058), .A0N(n2961), .A1N(n1722), .Y(n2968) );
  OAI211XL U2041 ( .A0(n3021), .A1(n1722), .B0(n1746), .C0(n3024), .Y(N665) );
  OAI211XL U2042 ( .A0(n2846), .A1(n1722), .B0(n2839), .C0(n2838), .Y(N721) );
  OAI211XL U2043 ( .A0(n3002), .A1(n1722), .B0(n3007), .C0(n3008), .Y(N679) );
  OAI211XL U2044 ( .A0(n3031), .A1(n1722), .B0(n3036), .C0(n3037), .Y(N651) );
  OAI211XL U2045 ( .A0(n1716), .A1(n3021), .B0(n1752), .C0(n3023), .Y(N666) );
  OAI211XL U2046 ( .A0(n1716), .A1(n2846), .B0(n2841), .C0(n2840), .Y(N722) );
  OAI211XL U2047 ( .A0(n1716), .A1(n3002), .B0(n3005), .C0(n3006), .Y(N680) );
  OAI211XL U2048 ( .A0(n3031), .A1(n1716), .B0(n3034), .C0(n3035), .Y(N652) );
  AOI22X2 U2049 ( .A0(n2366), .A1(n808), .B0(n2367), .B1(n807), .Y(n2369) );
  OAI211X2 U2050 ( .A0(n2366), .A1(n808), .B0(n2365), .C0(n809), .Y(n2370) );
  OAI211XL U2051 ( .A0(n1717), .A1(n3002), .B0(n3014), .C0(n3015), .Y(N675) );
  INVX3 U2052 ( .A(n1130), .Y(HC2[0]) );
  INVX3 U2053 ( .A(n1121), .Y(HC6[0]) );
  INVX3 U2054 ( .A(n1133), .Y(HC2[4]) );
  INVX3 U2055 ( .A(n1124), .Y(HC6[4]) );
  INVX3 U2056 ( .A(n1132), .Y(HC2[3]) );
  INVX3 U2057 ( .A(n1123), .Y(HC6[3]) );
  OAI211XL U2058 ( .A0(n1717), .A1(n3021), .B0(n1753), .C0(n3029), .Y(N661) );
  OAI211XL U2059 ( .A0(n1717), .A1(n2846), .B0(n2832), .C0(n2831), .Y(N717) );
  INVX3 U2060 ( .A(n1131), .Y(HC2[1]) );
  INVX3 U2061 ( .A(n1122), .Y(HC6[1]) );
  INVX3 U2062 ( .A(n1125), .Y(HC4[0]) );
  INVX3 U2063 ( .A(n1129), .Y(HC4[4]) );
  INVX3 U2064 ( .A(n1128), .Y(HC4[3]) );
  INVX3 U2065 ( .A(n1127), .Y(HC4[2]) );
  INVX3 U2066 ( .A(n1126), .Y(HC4[1]) );
  AOI22XL U2067 ( .A0(n1134), .A1(n3053), .B0(n2775), .B1(n3051), .Y(n3032) );
  AOI22XL U2068 ( .A0(n1134), .A1(n3056), .B0(n2775), .B1(n3054), .Y(n3034) );
  NAND2XL U2069 ( .A(n2775), .B(n3062), .Y(n2740) );
  AOI2BB2XL U2070 ( .B0(n2775), .B1(n3058), .A0N(n3038), .A1N(n1713), .Y(n3037) );
  AOI2BB2XL U2071 ( .B0(n2775), .B1(n3069), .A0N(n3038), .A1N(n1733), .Y(n3044) );
  NOR2XL U2072 ( .A(n1116), .B(n3021), .Y(n2791) );
  NOR2XL U2073 ( .A(n1116), .B(n3002), .Y(n2808) );
  NOR2XL U2074 ( .A(n1116), .B(n3031), .Y(n2774) );
  NOR2XL U2075 ( .A(n1116), .B(n2846), .Y(n2823) );
  CLKINVX1 U2077 ( .A(n2933), .Y(n1692) );
  OR2X1 U2078 ( .A(n2933), .B(n2349), .Y(n2644) );
  NOR2XL U2079 ( .A(n630), .B(n808), .Y(n2336) );
  OAI21XL U2080 ( .A0(n1864), .A1(n664), .B0(n1863), .Y(n850) );
  CLKINVX2 U2081 ( .A(n1251), .Y(n2801) );
  OAI211XL U2082 ( .A0(n2846), .A1(n1714), .B0(n2835), .C0(n2834), .Y(N716) );
  OAI211XL U2083 ( .A0(n3021), .A1(n1714), .B0(n1747), .C0(n3030), .Y(N660) );
  OAI211XL U2084 ( .A0(n3031), .A1(n1714), .B0(n3043), .C0(n3044), .Y(N646) );
  OAI211XL U2085 ( .A0(n3002), .A1(n1714), .B0(n3016), .C0(n3017), .Y(N674) );
  AOI22XL U2086 ( .A0(n1134), .A1(n3067), .B0(n2775), .B1(n3064), .Y(n3041) );
  NAND2XL U2087 ( .A(n2905), .B(n3064), .Y(n2974) );
  OAI211XL U2088 ( .A0(n1718), .A1(n2987), .B0(n1748), .C0(n2988), .Y(N695) );
  OAI211XL U2089 ( .A0(n1716), .A1(n2987), .B0(n1749), .C0(n2989), .Y(N694) );
  OAI211XL U2090 ( .A0(n1717), .A1(n2987), .B0(n1750), .C0(n2996), .Y(N689) );
  OAI211XL U2091 ( .A0(n2987), .A1(n1722), .B0(n1744), .C0(n2990), .Y(N693) );
  OAI211XL U2092 ( .A0(n2987), .A1(n1714), .B0(n1745), .C0(n2997), .Y(N688) );
  NOR2XL U2093 ( .A(n1116), .B(n2987), .Y(n2813) );
  OR2X2 U2094 ( .A(n2960), .B(n2677), .Y(n2987) );
  NAND3X4 U2095 ( .A(n2978), .B(n2961), .C(n2966), .Y(N700) );
  OAI211XL U2096 ( .A0(n1718), .A1(n2961), .B0(n2962), .C0(n2963), .Y(N709) );
  OAI211XL U2097 ( .A0(n1716), .A1(n2961), .B0(n2964), .C0(n2965), .Y(N708) );
  OAI211XL U2098 ( .A0(n1717), .A1(n2961), .B0(n2973), .C0(n2974), .Y(N703) );
  NOR2XL U2099 ( .A(n1116), .B(n2961), .Y(n2818) );
  NAND3X2 U2100 ( .A(n2733), .B(n2669), .C(n2982), .Y(n2961) );
  AOI21XL U2101 ( .A0(n2857), .A1(n3058), .B0(n2836), .Y(n2839) );
  AOI21XL U2102 ( .A0(n2857), .A1(n3069), .B0(n2833), .Y(n2835) );
  NAND2XL U2103 ( .A(n2857), .B(n3051), .Y(n2844) );
  NAND2XL U2104 ( .A(n2857), .B(n3054), .Y(n2840) );
  NOR2X2 U2105 ( .A(n2954), .B(n2653), .Y(n2857) );
  OAI21XL U2106 ( .A0(n1864), .A1(n671), .B0(n1862), .Y(n857) );
  OAI21XL U2107 ( .A0(n1875), .A1(n687), .B0(n1873), .Y(n873) );
  INVX3 U2108 ( .A(n2782), .Y(n2850) );
  INVX3 U2109 ( .A(n1086), .Y(n1794) );
  AOI2BB2XL U2110 ( .B0(n3064), .B1(n2583), .A0N(n2937), .A1N(n775), .Y(n2584)
         );
  NAND4X4 U2111 ( .A(n2749), .B(n3040), .C(n2848), .D(n2847), .Y(N644) );
  OAI21XL U2112 ( .A0(n1864), .A1(n670), .B0(n1861), .Y(n856) );
  OAI21XL U2113 ( .A0(n1864), .A1(n665), .B0(n1856), .Y(n851) );
  OAI21XL U2114 ( .A0(n1875), .A1(n681), .B0(n1867), .Y(n867) );
  OAI21XL U2115 ( .A0(n1875), .A1(n683), .B0(n1869), .Y(n869) );
  INVX4 U2116 ( .A(n1933), .Y(n1514) );
  NAND2X8 U2117 ( .A(n2246), .B(CNT6[6]), .Y(n2127) );
  AOI2BB2X4 U2118 ( .B0(n2049), .B1(n1976), .A0N(n1973), .A1N(n1758), .Y(n1366) );
  MXI2X4 U2119 ( .A(CNT4[5]), .B(n2001), .S0(n1786), .Y(n1758) );
  NAND2X8 U2120 ( .A(n1578), .B(n1644), .Y(n2156) );
  INVX8 U2121 ( .A(n2295), .Y(n2209) );
  NAND2X4 U2122 ( .A(n2296), .B(n2209), .Y(n2193) );
  NAND2X6 U2123 ( .A(n1406), .B(n1373), .Y(n1401) );
  AND2X8 U2124 ( .A(n1959), .B(n1269), .Y(n1687) );
  NAND2X2 U2125 ( .A(n1941), .B(n1943), .Y(n1270) );
  INVX8 U2126 ( .A(n1557), .Y(n1755) );
  NAND2X4 U2127 ( .A(n2242), .B(n2421), .Y(n2243) );
  NAND2X8 U2128 ( .A(n1272), .B(n1069), .Y(n2101) );
  NAND2X8 U2129 ( .A(n2036), .B(n2037), .Y(n1624) );
  NAND2X8 U2130 ( .A(n2214), .B(n2287), .Y(n2196) );
  MXI2X4 U2131 ( .A(n1329), .B(CNT5[5]), .S0(n1690), .Y(n1338) );
  MXI2X2 U2132 ( .A(n1000), .B(n1977), .S0(n1339), .Y(n2090) );
  AOI21X4 U2133 ( .A0(n2067), .A1(n2066), .B0(n1481), .Y(n1375) );
  AND2X8 U2134 ( .A(n1276), .B(n1959), .Y(n1689) );
  INVX12 U2135 ( .A(n1935), .Y(n1972) );
  CLKAND2X12 U2136 ( .A(n2094), .B(n1979), .Y(n1990) );
  NAND2X6 U2137 ( .A(n1984), .B(n1950), .Y(n1675) );
  AND3X8 U2138 ( .A(n1277), .B(n2101), .C(n2100), .Y(n1643) );
  BUFX4 U2139 ( .A(n2078), .Y(n1278) );
  AND2X8 U2140 ( .A(n1578), .B(n1645), .Y(n1575) );
  NAND2X6 U2141 ( .A(n2200), .B(n2192), .Y(n1282) );
  NAND2X6 U2142 ( .A(n1566), .B(n2104), .Y(n2105) );
  NAND2X8 U2143 ( .A(n1637), .B(n2256), .Y(n1634) );
  NAND2X6 U2144 ( .A(n1390), .B(n1388), .Y(n1387) );
  OAI22X4 U2145 ( .A0(n1568), .A1(n1567), .B0(n1763), .B1(n2415), .Y(n2098) );
  NOR2X8 U2146 ( .A(n1773), .B(n2213), .Y(n2102) );
  NAND2X4 U2147 ( .A(n2409), .B(n2230), .Y(n2211) );
  NOR2X8 U2148 ( .A(n1680), .B(n1689), .Y(n1359) );
  NAND3X8 U2149 ( .A(n1365), .B(n1681), .C(n1364), .Y(n1363) );
  NAND3X8 U2150 ( .A(n1363), .B(n1361), .C(n1362), .Y(n1963) );
  AND2X8 U2151 ( .A(n2016), .B(n1289), .Y(n2027) );
  MXI2X4 U2152 ( .A(n1514), .B(n1018), .S0(n1217), .Y(n1968) );
  OR2X8 U2153 ( .A(n1384), .B(n954), .Y(n1636) );
  MXI2X4 U2154 ( .A(n947), .B(n1760), .S0(n1494), .Y(n1319) );
  MXI2X4 U2155 ( .A(n1218), .B(n2150), .S0(n1648), .Y(n2270) );
  NAND2X6 U2156 ( .A(n2223), .B(n2410), .Y(n2238) );
  NAND2X8 U2157 ( .A(n2289), .B(n2191), .Y(n2192) );
  INVX16 U2158 ( .A(n2127), .Y(n2128) );
  NAND2X6 U2159 ( .A(n2193), .B(n2199), .Y(n1281) );
  BUFX4 U2160 ( .A(n1772), .Y(n1283) );
  MXI2X4 U2161 ( .A(n1761), .B(n2289), .S0(n982), .Y(n2230) );
  NOR2X8 U2162 ( .A(n1538), .B(n1537), .Y(n1536) );
  CLKBUFX3 U2163 ( .A(n2395), .Y(n1285) );
  NOR2X8 U2164 ( .A(n2254), .B(n2255), .Y(n2160) );
  NOR2X8 U2165 ( .A(n1286), .B(n2201), .Y(n1662) );
  NOR2X8 U2166 ( .A(n1759), .B(n2399), .Y(n1566) );
  INVX6 U2167 ( .A(n2190), .Y(n2289) );
  AND3X8 U2168 ( .A(n2154), .B(n2155), .C(n2159), .Y(n1776) );
  AND2X8 U2169 ( .A(n1914), .B(n1614), .Y(n1295) );
  NOR2X6 U2170 ( .A(n2067), .B(n2066), .Y(n1417) );
  INVX12 U2171 ( .A(n1422), .Y(n1799) );
  NAND2X8 U2172 ( .A(n1604), .B(n1105), .Y(n1287) );
  NAND2X4 U2173 ( .A(n2055), .B(n2134), .Y(n2053) );
  NAND2X6 U2174 ( .A(n2128), .B(CNT6[7]), .Y(n2129) );
  MXI2X4 U2175 ( .A(n2115), .B(n671), .S0(n1690), .Y(n2151) );
  BUFX4 U2176 ( .A(n2418), .Y(n1291) );
  NAND2BX2 U2177 ( .AN(n605), .B(n2592), .Y(n2593) );
  NAND2BX2 U2178 ( .AN(n606), .B(n2592), .Y(n2590) );
  AND2X8 U2179 ( .A(n2231), .B(n2211), .Y(n2241) );
  BUFX4 U2180 ( .A(n2052), .Y(n1294) );
  INVX6 U2181 ( .A(n1987), .Y(n2087) );
  NAND2X4 U2182 ( .A(n2415), .B(n1763), .Y(n1542) );
  OA21X4 U2183 ( .A0(n2259), .A1(n2181), .B0(n2149), .Y(n1724) );
  NAND3X8 U2184 ( .A(n1109), .B(n1724), .C(n1576), .Y(n2158) );
  INVX8 U2185 ( .A(n2219), .Y(n2220) );
  NAND2X6 U2186 ( .A(n2297), .B(n2298), .Y(n2194) );
  INVX3 U2187 ( .A(n1293), .Y(n2212) );
  NAND2BX4 U2188 ( .AN(n1215), .B(n1525), .Y(n1955) );
  INVX4 U2189 ( .A(n1663), .Y(n1661) );
  NAND2X6 U2190 ( .A(n2032), .B(CNT5[7]), .Y(n2033) );
  NAND3X6 U2191 ( .A(n1378), .B(n1380), .C(n1377), .Y(n1376) );
  NAND2X6 U2192 ( .A(n1630), .B(n1297), .Y(n1423) );
  NOR2X8 U2193 ( .A(n1298), .B(n1299), .Y(n1297) );
  NAND2X8 U2194 ( .A(n2195), .B(n2201), .Y(n1298) );
  MXI2X4 U2195 ( .A(n2007), .B(n679), .S0(n1786), .Y(n2040) );
  NAND2X2 U2196 ( .A(n2040), .B(n671), .Y(n2008) );
  CLKBUFX3 U2197 ( .A(n2188), .Y(n1301) );
  MXI2X8 U2198 ( .A(n2087), .B(n1317), .S0(n1499), .Y(n1762) );
  OAI21X4 U2199 ( .A0(n2091), .A1(n1492), .B0(n1303), .Y(n1407) );
  AOI22X2 U2200 ( .A0(n630), .A1(\com[2][1] ), .B0(\com[2][2] ), .B1(n631), 
        .Y(n2306) );
  NAND2X2 U2201 ( .A(n1773), .B(n2213), .Y(n2099) );
  NAND2BX4 U2202 ( .AN(n2603), .B(n2417), .Y(n1309) );
  NOR2X8 U2203 ( .A(n2004), .B(n2005), .Y(n2012) );
  NAND2X4 U2204 ( .A(n2401), .B(n1307), .Y(n1306) );
  NAND2X6 U2205 ( .A(n2450), .B(n2595), .Y(n2433) );
  BUFX4 U2206 ( .A(n2613), .Y(n1308) );
  NAND2X8 U2207 ( .A(n1420), .B(n1772), .Y(n2236) );
  INVXL U2208 ( .A(n2136), .Y(n1686) );
  BUFX4 U2209 ( .A(n2255), .Y(n1312) );
  BUFX20 U2210 ( .A(n2385), .Y(n1773) );
  BUFX4 U2211 ( .A(n2406), .Y(n1314) );
  NAND2X8 U2212 ( .A(n1315), .B(n1622), .Y(n1605) );
  MXI2X6 U2213 ( .A(n1971), .B(n1972), .S0(n1787), .Y(n1970) );
  NAND2BX2 U2214 ( .AN(n607), .B(n2592), .Y(n2589) );
  NAND2X8 U2215 ( .A(n1605), .B(n1600), .Y(n1355) );
  NAND2X6 U2216 ( .A(n2080), .B(n2068), .Y(n1373) );
  NOR2X8 U2217 ( .A(n1316), .B(n1355), .Y(n1357) );
  INVX12 U2218 ( .A(n1397), .Y(n1949) );
  MXI2X8 U2219 ( .A(n2174), .B(n955), .S0(n1383), .Y(n2298) );
  OA21X4 U2220 ( .A0(n2070), .A1(n2139), .B0(n1310), .Y(n1372) );
  AOI21X4 U2221 ( .A0(n1470), .A1(n1469), .B0(n1320), .Y(n1468) );
  BUFX4 U2222 ( .A(n2410), .Y(n1322) );
  OAI21X4 U2223 ( .A0(n1947), .A1(n1092), .B0(n1512), .Y(n1511) );
  INVX6 U2224 ( .A(n2141), .Y(n2246) );
  OAI2BB1X4 U2225 ( .A0N(CNT4[4]), .A1N(n1917), .B0(n1328), .Y(n1623) );
  NAND2X4 U2226 ( .A(n1952), .B(CNT4[3]), .Y(n1328) );
  NAND2X2 U2227 ( .A(n1319), .B(n1756), .Y(n2185) );
  INVX12 U2228 ( .A(n2614), .Y(n2623) );
  NOR2X8 U2229 ( .A(n1333), .B(n1507), .Y(n1503) );
  NAND2X8 U2230 ( .A(n1657), .B(n1656), .Y(n1335) );
  MXI2X4 U2231 ( .A(n1198), .B(n1238), .S0(n1343), .Y(n1500) );
  OAI2BB1X4 U2233 ( .A0N(n1345), .A1N(n2769), .B0(n1344), .Y(n2772) );
  NAND2X8 U2234 ( .A(n1348), .B(n1587), .Y(n1347) );
  OAI2BB1X4 U2235 ( .A0N(n1931), .A1N(n1353), .B0(n1354), .Y(n1973) );
  MXI2X4 U2236 ( .A(n1977), .B(n1000), .S0(n1787), .Y(n1976) );
  INVX20 U2237 ( .A(n1357), .Y(n1786) );
  NAND2X8 U2238 ( .A(n1358), .B(n1683), .Y(n1962) );
  NOR2X8 U2239 ( .A(n1688), .B(n1689), .Y(n1361) );
  OR2X8 U2240 ( .A(n2097), .B(n1988), .Y(n1993) );
  AOI21X4 U2241 ( .A0(n2064), .A1(n1419), .B0(n1370), .Y(n1369) );
  OAI21X4 U2242 ( .A0(n2054), .A1(n2150), .B0(n2053), .Y(n1371) );
  NAND2X4 U2243 ( .A(n2135), .B(n1379), .Y(n1418) );
  MXI2X4 U2244 ( .A(n2041), .B(n2042), .S0(n1673), .Y(n2080) );
  OR2X8 U2245 ( .A(n2069), .B(n2081), .Y(n1406) );
  MXI2X4 U2246 ( .A(n1004), .B(n1294), .S0(n1367), .Y(n2069) );
  MXI2X4 U2247 ( .A(n1493), .B(n2049), .S0(n1646), .Y(n2060) );
  MXI2X4 U2248 ( .A(n1294), .B(n1004), .S0(n1374), .Y(n2134) );
  MXI2X4 U2249 ( .A(n2049), .B(n1493), .S0(n1374), .Y(n2091) );
  NAND2X4 U2250 ( .A(n1473), .B(n2086), .Y(n1524) );
  NAND2X8 U2251 ( .A(n2435), .B(n2613), .Y(n1381) );
  NAND3X6 U2252 ( .A(n1382), .B(n1442), .C(n1435), .Y(n1441) );
  NAND3X6 U2253 ( .A(n1382), .B(n1442), .C(n1439), .Y(n1438) );
  NAND3X8 U2254 ( .A(n1503), .B(n1502), .C(n1504), .Y(n1382) );
  NAND2X8 U2255 ( .A(n1555), .B(n1384), .Y(n2576) );
  NAND2X8 U2256 ( .A(n1430), .B(n1429), .Y(n1384) );
  NAND3X6 U2257 ( .A(n1384), .B(n1574), .C(n1572), .Y(n1635) );
  NOR2X6 U2258 ( .A(n2153), .B(n1556), .Y(n1386) );
  NAND2BX4 U2259 ( .AN(n1651), .B(n1389), .Y(n1388) );
  AND2X8 U2260 ( .A(n2161), .B(n2252), .Y(n1652) );
  AND2X8 U2261 ( .A(n1571), .B(n2251), .Y(n1651) );
  MXI2X4 U2262 ( .A(n1216), .B(n2135), .S0(n1195), .Y(n2144) );
  MXI2X4 U2263 ( .A(n1085), .B(n2133), .S0(n1195), .Y(n2165) );
  MXI2X4 U2264 ( .A(n1771), .B(n1431), .S0(n1195), .Y(n2263) );
  NOR2X6 U2265 ( .A(n1395), .B(n1394), .Y(n1393) );
  NAND2X4 U2266 ( .A(n2122), .B(n2121), .Y(n1395) );
  NAND2X4 U2267 ( .A(n2141), .B(n681), .Y(n2121) );
  NAND3X6 U2268 ( .A(n1093), .B(n1528), .C(n1106), .Y(n2126) );
  INVX6 U2269 ( .A(n1396), .Y(n2188) );
  CLKMX2X6 U2270 ( .A(n1916), .B(n657), .S0(n1137), .Y(n1397) );
  MXI2X4 U2271 ( .A(n2039), .B(n2038), .S0(n981), .Y(n2131) );
  MXI2X4 U2272 ( .A(n1408), .B(n1003), .S0(n1494), .Y(n2385) );
  NAND2BX4 U2273 ( .AN(n2445), .B(n2597), .Y(n1669) );
  MXI2X4 U2274 ( .A(n1413), .B(n999), .S0(n930), .Y(n2445) );
  NAND3X2 U2275 ( .A(n2425), .B(n1414), .C(n2623), .Y(n2420) );
  NAND2X6 U2276 ( .A(n1410), .B(n1672), .Y(n1415) );
  NAND2X6 U2277 ( .A(n2596), .B(n2451), .Y(n2432) );
  MXI2X4 U2278 ( .A(n2212), .B(n2213), .S0(n1638), .Y(n2224) );
  OR2X8 U2279 ( .A(n1651), .B(n1652), .Y(n1429) );
  AND2X8 U2280 ( .A(n1518), .B(n1918), .Y(n1432) );
  OR2X8 U2281 ( .A(n1919), .B(n1434), .Y(n1433) );
  MXI2X8 U2282 ( .A(CNT1[5]), .B(CNT2[5]), .S0(n1784), .Y(n1609) );
  AND2X8 U2283 ( .A(n1915), .B(CNT4[5]), .Y(n1919) );
  AND2X8 U2284 ( .A(n1768), .B(n1236), .Y(n1893) );
  NAND3X8 U2285 ( .A(n1908), .B(n1906), .C(n1907), .Y(n1442) );
  NAND2X8 U2286 ( .A(n1438), .B(n1621), .Y(n1437) );
  AOI2BB1X4 U2287 ( .A0N(n1909), .A1N(n656), .B0(n1500), .Y(n1440) );
  NOR2X6 U2288 ( .A(n1770), .B(n1212), .Y(n1887) );
  OAI21X4 U2289 ( .A0(n1885), .A1(n1206), .B0(n1884), .Y(n1890) );
  MXI2X4 U2292 ( .A(n2600), .B(n2598), .S0(n1803), .Y(\com[4][1] ) );
  NAND2BX4 U2302 ( .AN(n2629), .B(n608), .Y(n1460) );
  MXI2X4 U2303 ( .A(n1308), .B(n2612), .S0(n1352), .Y(n2630) );
  MXI2X4 U2307 ( .A(n2434), .B(n2611), .S0(n1352), .Y(n1464) );
  MXI2X4 U2309 ( .A(n2615), .B(n2614), .S0(n1352), .Y(n1466) );
  NAND2X4 U2310 ( .A(n2299), .B(n1468), .Y(n2303) );
  OAI22X4 U2311 ( .A0(\com[3][0] ), .A1(n629), .B0(n630), .B1(\com[3][1] ), 
        .Y(n1469) );
  OAI21X4 U2312 ( .A0(n979), .A1(n2279), .B0(n1522), .Y(\com[3][0] ) );
  AOI22X4 U2313 ( .A0(\com[3][1] ), .A1(n630), .B0(n1100), .B1(n631), .Y(n1470) );
  CLKMX2X6 U2314 ( .A(n2387), .B(n1247), .S0(n1313), .Y(n1467) );
  OAI2BB2X4 U2315 ( .B0(n1288), .B1(n1472), .A0N(n2091), .A1N(n1492), .Y(n1471) );
  CLKINVX6 U2316 ( .A(n2087), .Y(n1472) );
  MXI2X4 U2317 ( .A(n2268), .B(n2170), .S0(n1193), .Y(n2291) );
  MXI2X4 U2318 ( .A(n1002), .B(n1177), .S0(n1646), .Y(n1980) );
  MXI2X4 U2319 ( .A(n2182), .B(n2181), .S0(n1474), .Y(n2288) );
  NAND2X8 U2320 ( .A(n1005), .B(n1962), .Y(n1646) );
  INVX8 U2321 ( .A(n1761), .Y(n2191) );
  OAI2BB1X4 U2322 ( .A0N(CNT5[3]), .A1N(n2045), .B0(n1289), .Y(n2004) );
  NAND4X8 U2323 ( .A(n1536), .B(n1535), .C(n1534), .D(n1542), .Y(n1642) );
  NAND2X2 U2324 ( .A(n1947), .B(n1092), .Y(n1924) );
  NAND2X4 U2325 ( .A(n1761), .B(n2190), .Y(n2197) );
  INVX8 U2326 ( .A(n2406), .Y(n1568) );
  INVX4 U2327 ( .A(n2425), .Y(n2423) );
  INVX20 U2328 ( .A(n1519), .Y(n1582) );
  INVX6 U2330 ( .A(n1973), .Y(n2048) );
  NAND2X6 U2331 ( .A(n1592), .B(n1593), .Y(n1603) );
  NAND2X4 U2332 ( .A(n2601), .B(n2447), .Y(n2396) );
  NOR2X8 U2333 ( .A(n1619), .B(n2077), .Y(n2078) );
  NAND3X8 U2334 ( .A(n1636), .B(n1635), .C(n1634), .Y(n1691) );
  MXI2X4 U2335 ( .A(n1225), .B(n670), .S0(n1690), .Y(n2114) );
  AOI22X2 U2336 ( .A0(n686), .A1(n2114), .B0(n2151), .B1(n687), .Y(n1529) );
  NAND2X8 U2338 ( .A(n2180), .B(n2085), .Y(n1627) );
  MXI2X1 U2339 ( .A(n2598), .B(n2600), .S0(n1352), .Y(n2608) );
  MXI2X4 U2340 ( .A(n677), .B(n1332), .S0(n1786), .Y(n2049) );
  MXI2X4 U2341 ( .A(n1966), .B(n968), .S0(n1217), .Y(n2042) );
  NAND2X8 U2342 ( .A(n2138), .B(n2137), .Y(n2152) );
  NAND2BX4 U2343 ( .AN(n2060), .B(n1045), .Y(n1478) );
  NAND2X4 U2344 ( .A(n2285), .B(n1565), .Y(n2421) );
  MXI2X4 U2345 ( .A(n2075), .B(n2077), .S0(n1076), .Y(n2285) );
  NOR2X6 U2350 ( .A(\com[4][6] ), .B(n1112), .Y(n1486) );
  NAND2X4 U2351 ( .A(n1489), .B(n2454), .Y(n1488) );
  NAND2X4 U2352 ( .A(\com[4][6] ), .B(n614), .Y(n1489) );
  BUFX20 U2354 ( .A(n1075), .Y(n1494) );
  NAND3X8 U2355 ( .A(n1497), .B(n1495), .C(n1496), .Y(n1659) );
  NAND3X8 U2356 ( .A(n1545), .B(n1546), .C(n1585), .Y(n1495) );
  MXI2X4 U2357 ( .A(n1085), .B(n2133), .S0(n1791), .Y(n2267) );
  OAI21X4 U2358 ( .A0(n2268), .A1(n2270), .B0(n1498), .Y(n1576) );
  MXI2X4 U2359 ( .A(CNT6[1]), .B(n2114), .S0(n1569), .Y(n2266) );
  MXI2X4 U2360 ( .A(n1015), .B(n2258), .S0(n2576), .Y(n2215) );
  CLKAND2X12 U2361 ( .A(n1508), .B(n1509), .Y(n1908) );
  MXI2X4 U2362 ( .A(n1926), .B(n1925), .S0(n1024), .Y(n1969) );
  OAI2BB1X4 U2363 ( .A0N(n1953), .A1N(n1967), .B0(n1924), .Y(n1516) );
  MXI2X4 U2364 ( .A(CNT3[0]), .B(n1923), .S0(n1326), .Y(n1967) );
  CLKMX2X6 U2365 ( .A(n1927), .B(CNT3[3]), .S0(n1137), .Y(n1517) );
  AND3X8 U2366 ( .A(n1518), .B(n1918), .C(CNT4[7]), .Y(n1611) );
  MXI2X4 U2367 ( .A(n1010), .B(n1520), .S0(n1799), .Y(n1521) );
  MXI2X4 U2368 ( .A(n2291), .B(n1523), .S0(n1331), .Y(\com[2][0] ) );
  MXI2X4 U2369 ( .A(n1267), .B(n2286), .S0(n1331), .Y(\com[2][6] ) );
  MXI2X4 U2370 ( .A(n1527), .B(n1988), .S0(n1582), .Y(n1557) );
  MXI2X4 U2371 ( .A(n1997), .B(n1998), .S0(n1526), .Y(n2075) );
  MXI2X4 U2372 ( .A(n2081), .B(n2082), .S0(n1526), .Y(n2390) );
  MXI2X4 U2373 ( .A(n2087), .B(n1317), .S0(n1526), .Y(n2415) );
  AOI2BB1X4 U2374 ( .A0N(n2118), .A1N(n685), .B0(n1529), .Y(n1528) );
  NAND3X6 U2375 ( .A(n2124), .B(n2125), .C(n1082), .Y(n1532) );
  OAI2BB1X4 U2376 ( .A0N(n684), .A1N(n2120), .B0(n2119), .Y(n2124) );
  NAND3X6 U2377 ( .A(n1642), .B(n1641), .C(n1640), .Y(n1558) );
  MXI2X4 U2378 ( .A(n2083), .B(n949), .S0(n1793), .Y(n2389) );
  NAND2X6 U2379 ( .A(n2395), .B(n2203), .Y(n1541) );
  MXI2X4 U2380 ( .A(n2163), .B(n2162), .S0(n1193), .Y(n2293) );
  NAND2X8 U2381 ( .A(n1633), .B(n1547), .Y(n1546) );
  NOR2X8 U2382 ( .A(n2153), .B(n1556), .Y(n1650) );
  INVX12 U2383 ( .A(n1651), .Y(n1556) );
  NAND3X6 U2384 ( .A(n1642), .B(n1643), .C(n1641), .Y(n1559) );
  NAND2X8 U2385 ( .A(n1560), .B(n1570), .Y(n2138) );
  NAND2X8 U2386 ( .A(n1562), .B(n1561), .Y(n2137) );
  AND2X8 U2387 ( .A(n2129), .B(n2130), .Y(n1561) );
  NOR2X8 U2388 ( .A(n2285), .B(n1564), .Y(n1663) );
  MXI2X4 U2389 ( .A(n950), .B(n2089), .S0(n1792), .Y(n2406) );
  AND2X8 U2390 ( .A(n2127), .B(n680), .Y(n1570) );
  MXI2X4 U2391 ( .A(CNT6[6]), .B(n2141), .S0(n2152), .Y(n2255) );
  MXI2X4 U2392 ( .A(n1222), .B(n2167), .S0(n1076), .Y(n2395) );
  ACHCINX2 U2393 ( .CIN(n1580), .A(n2165), .B(n2164), .CO(n1585) );
  AOI2BB2X4 U2394 ( .B0(n1582), .B1(n2081), .A0N(n1582), .A1N(n1579), .Y(n2164) );
  NAND2X4 U2395 ( .A(n2167), .B(n2168), .Y(n1580) );
  AOI2BB2X4 U2396 ( .B0(n1582), .B1(n2079), .A0N(n1582), .A1N(n1581), .Y(n2167) );
  MXI2X4 U2397 ( .A(n1203), .B(n1214), .S0(n1784), .Y(n1923) );
  OAI21X4 U2398 ( .A0(n1245), .A1(n1880), .B0(n1879), .Y(n1589) );
  AOI22X4 U2399 ( .A0(n1999), .A1(n1618), .B0(n672), .B1(n673), .Y(n1592) );
  OAI21X4 U2400 ( .A0(n1999), .A1(n672), .B0(n1949), .Y(n1593) );
  AND2X8 U2401 ( .A(n1942), .B(n1946), .Y(n1594) );
  NAND3X6 U2402 ( .A(n1940), .B(n1596), .C(n1597), .Y(n1595) );
  AOI2BB1X4 U2403 ( .A0N(n1513), .A1N(n1937), .B0(n1598), .Y(n1597) );
  NAND2X4 U2404 ( .A(n1933), .B(n1969), .Y(n1937) );
  NAND3X6 U2405 ( .A(n1601), .B(n1603), .C(n1920), .Y(n1600) );
  AOI22X4 U2406 ( .A0(n2002), .A1(n676), .B0(n2009), .B1(n677), .Y(n1602) );
  NAND3X6 U2407 ( .A(n1940), .B(n1607), .C(n1596), .Y(n1936) );
  NOR2X6 U2408 ( .A(n1608), .B(n1674), .Y(n1607) );
  OAI21X4 U2409 ( .A0(n2000), .A1(CNT4[1]), .B0(n1613), .Y(n1612) );
  NAND2X4 U2410 ( .A(n2006), .B(n679), .Y(n1613) );
  MXI2X4 U2411 ( .A(n1912), .B(n663), .S0(n1024), .Y(n2006) );
  AOI22X4 U2412 ( .A0(n2000), .A1(CNT4[1]), .B0(n1952), .B1(CNT4[3]), .Y(n1614) );
  MXI2X4 U2413 ( .A(n1615), .B(CNT3[1]), .S0(n1025), .Y(n2000) );
  AOI22X4 U2414 ( .A0(CNT4[5]), .A1(n1915), .B0(CNT4[4]), .B1(n1917), .Y(n1616) );
  NAND2X4 U2415 ( .A(n1971), .B(n1935), .Y(n1617) );
  NAND2BX4 U2416 ( .AN(n672), .B(CNT4[6]), .Y(n1618) );
  INVX1 U2417 ( .A(n1949), .Y(n2014) );
  AND2X6 U2418 ( .A(n1909), .B(n656), .Y(n1621) );
  AND2X8 U2419 ( .A(n2076), .B(n2077), .Y(n1628) );
  OR2X8 U2420 ( .A(n2198), .B(n2197), .Y(n1630) );
  CLKINVX20 U2421 ( .A(n1638), .Y(n1639) );
  MXI2X4 U2422 ( .A(n684), .B(n2248), .S0(n2152), .Y(n2261) );
  NAND2X6 U2423 ( .A(n2261), .B(n2263), .Y(n1645) );
  OAI21X4 U2424 ( .A0(n2261), .A1(n2263), .B0(n2146), .Y(n1647) );
  NAND2X8 U2425 ( .A(n2255), .B(n2254), .Y(n2154) );
  NAND2X4 U2426 ( .A(n2144), .B(n2257), .Y(n2155) );
  AND2X8 U2427 ( .A(n1993), .B(n1997), .Y(n1654) );
  MXI2X4 U2428 ( .A(n1337), .B(n2166), .S0(n1792), .Y(n2292) );
  NOR2BX4 U2429 ( .AN(n2308), .B(n1664), .Y(n2480) );
  NAND2X4 U2430 ( .A(\com[2][5] ), .B(n634), .Y(n2311) );
  MXI2X4 U2431 ( .A(n2295), .B(n2296), .S0(n1331), .Y(\com[2][3] ) );
  NOR2X6 U2432 ( .A(n1666), .B(n1098), .Y(n1665) );
  NOR2X6 U2433 ( .A(n1667), .B(n2614), .Y(n1666) );
  NAND2X4 U2434 ( .A(n1675), .B(n1943), .Y(n1674) );
  OR2X8 U2435 ( .A(n1280), .B(CNT5[3]), .Y(n1677) );
  NAND2X4 U2436 ( .A(n1957), .B(n1958), .Y(n1680) );
  OAI2BB1X4 U2437 ( .A0N(n2042), .A1N(n1965), .B0(n1682), .Y(n1681) );
  AND2X6 U2438 ( .A(n2031), .B(n664), .Y(n1684) );
  INVX3 U2440 ( .A(n1100), .Y(n2367) );
  CLKINVX2 U2441 ( .A(n1639), .Y(n1795) );
  OAI21X4 U2442 ( .A0(n1420), .A1(n1772), .B0(n2218), .Y(n2219) );
  NAND2X2 U2443 ( .A(n2267), .B(n2163), .Y(n2148) );
  MXI2X4 U2444 ( .A(n2169), .B(n1223), .S0(n1076), .Y(n2290) );
  OAI21X4 U2445 ( .A0(n2051), .A1(n670), .B0(n2025), .Y(n2005) );
  MXI2X4 U2446 ( .A(n2150), .B(n1218), .S0(n1791), .Y(n2168) );
  OAI21X4 U2447 ( .A0(n2110), .A1(CNT5[1]), .B0(n2008), .Y(n2011) );
  MXI2X4 U2448 ( .A(CNT5[1]), .B(n1268), .S0(n1789), .Y(n2055) );
  AOI21X4 U2449 ( .A0(n2024), .A1(n1271), .B0(n2015), .Y(n2019) );
  NAND2X6 U2450 ( .A(n2173), .B(n2264), .Y(n2146) );
  NAND2X2 U2451 ( .A(n2045), .B(CNT5[3]), .Y(n2016) );
  AOI21X4 U2452 ( .A0(n2024), .A1(n1271), .B0(n2023), .Y(n2029) );
  NAND2X4 U2453 ( .A(n2225), .B(n2399), .Y(n2100) );
  NAND2X8 U2454 ( .A(n2111), .B(n666), .Y(n2022) );
  INVX8 U2455 ( .A(n2144), .Y(n2258) );
  MXI2X4 U2456 ( .A(n2180), .B(n945), .S0(n1076), .Y(n2190) );
  OAI22X2 U2458 ( .A0(n630), .A1(\com[2][1] ), .B0(\com[2][0] ), .B1(n629), 
        .Y(n2305) );
  MXI2X4 U2459 ( .A(n2209), .B(n2208), .S0(n982), .Y(n2414) );
  NAND2X2 U2460 ( .A(n2290), .B(n2291), .Y(n2176) );
  MXI2X1 U2461 ( .A(n1285), .B(n2394), .S0(n1796), .Y(n2447) );
  OA21X4 U2462 ( .A0(n2292), .A1(n2293), .B0(n2185), .Y(n1778) );
  CLKINVX8 U2463 ( .A(n2174), .Y(n2264) );
  NAND2X6 U2464 ( .A(n1757), .B(n1267), .Y(n2195) );
  NAND3X8 U2465 ( .A(n2012), .B(n2011), .C(n2010), .Y(n2030) );
  NAND2X2 U2466 ( .A(n2275), .B(n2405), .Y(n2232) );
  INVX3 U2468 ( .A(\com[3][4] ), .Y(n2372) );
  OAI22X1 U2469 ( .A0(n2357), .A1(\com[3][4] ), .B0(\com[3][3] ), .B1(n2356), 
        .Y(n2358) );
  OA21X4 U2470 ( .A0(n2414), .A1(n2233), .B0(n2211), .Y(n1710) );
  OAI2BB1X4 U2472 ( .A0N(n2233), .A1N(n2414), .B0(n2232), .Y(n2240) );
  OAI2BB1X4 U2475 ( .A0N(n668), .A1N(n2112), .B0(n2017), .Y(n2026) );
  CLKAND2X12 U2476 ( .A(n2222), .B(n2386), .Y(n1779) );
  OAI22X2 U2477 ( .A0(n2374), .A1(n2373), .B0(n2372), .B1(n805), .Y(n2375) );
  AO21X4 U2478 ( .A0(n1352), .A1(n2606), .B0(n2605), .Y(n2607) );
  OAI21X2 U2479 ( .A0(n623), .A1(\com[3][5] ), .B0(n2375), .Y(n2377) );
  OAI211X2 U2480 ( .A0(n3234), .A1(n3233), .B0(n2490), .C0(n3232), .Y(n776) );
  OAI2BB1X4 U2482 ( .A0N(n2295), .A1N(n2208), .B0(n2194), .Y(n2200) );
  OAI2BB1X4 U2484 ( .A0N(n1398), .A1N(n2047), .B0(n1956), .Y(n1960) );
  AOI21X2 U2486 ( .A0(n2370), .A1(n2369), .B0(n2368), .Y(n2374) );
  NAND2X4 U2487 ( .A(n1801), .B(n2419), .Y(n2425) );
  AOI21X4 U2488 ( .A0(n2177), .A1(n2176), .B0(n2175), .Y(n2187) );
  MXI2X4 U2489 ( .A(n1247), .B(n2387), .S0(n930), .Y(n2603) );
  MXI2X4 U2490 ( .A(n1540), .B(n1292), .S0(n1639), .Y(n2216) );
  INVX3 U2491 ( .A(\com[3][1] ), .Y(n2366) );
  MXI2X2 U2492 ( .A(n959), .B(n1983), .S0(n1339), .Y(n1988) );
  MXI2X1 U2493 ( .A(n1972), .B(n1971), .S0(n1339), .Y(n1987) );
  OAI211XL U2494 ( .A0(re_order_en), .A1(n3046), .B0(n2927), .C0(n2944), .Y(
        N204) );
  MXI2X1 U2495 ( .A(n2562), .B(n2561), .S0(n1780), .Y(n2573) );
  AOI211X1 U2496 ( .A0(tree_mem[1]), .A1(tree_mem[2]), .B0(tree_mem[0]), .C0(
        n2923), .Y(n2922) );
  NOR4X1 U2497 ( .A(tree_mem[0]), .B(tree_mem[1]), .C(n2923), .D(n1702), .Y(
        n2920) );
  NOR2X1 U2498 ( .A(n1712), .B(n3046), .Y(n2925) );
  XOR2X1 U2499 ( .A(n2928), .B(tree_mem_back[0]), .Y(n785) );
  OAI211X1 U2500 ( .A0(tree_mem_back[1]), .A1(n3069), .B0(n2939), .C0(n2473), 
        .Y(n2940) );
  AOI2BB2XL U2512 ( .B0(n2947), .B1(n533), .A0N(n2947), .A1N(n3085), .Y(n731)
         );
  AOI2BB2XL U2513 ( .B0(n2947), .B1(n535), .A0N(n2947), .A1N(n3080), .Y(n732)
         );
  AOI2BB2XL U2514 ( .B0(n2947), .B1(n540), .A0N(n1814), .A1N(n3094), .Y(n735)
         );
  AOI2BB2XL U2515 ( .B0(n2947), .B1(n538), .A0N(n1814), .A1N(n3099), .Y(n734)
         );
  AOI2BB2XL U2516 ( .B0(n2947), .B1(n531), .A0N(n1814), .A1N(n3095), .Y(n730)
         );
  BUFX12 U2517 ( .A(n2947), .Y(n1814) );
  NAND3X2 U2518 ( .A(state[2]), .B(state[0]), .C(n1725), .Y(n2947) );
  OAI2BB1X1 U2519 ( .A0N(n2284), .A1N(N1143), .B0(n2281), .Y(n814) );
  OAI2BB1X1 U2520 ( .A0N(n2284), .A1N(N1144), .B0(n2280), .Y(n815) );
  OAI2BB1X1 U2521 ( .A0N(n2284), .A1N(N1145), .B0(n2274), .Y(n816) );
  OAI2BB1X2 U2522 ( .A0N(n2284), .A1N(N1146), .B0(n2272), .Y(n817) );
  INVX3 U2524 ( .A(n2282), .Y(n2284) );
  NOR2X1 U2525 ( .A(n3109), .B(n3110), .Y(n2912) );
  CLKINVX1 U2526 ( .A(n2322), .Y(n2271) );
  CLKMX2X2 U2529 ( .A(n2772), .B(n3049), .S0(n2910), .Y(n770) );
  OAI21X1 U2530 ( .A0(n2768), .A1(\com[1][6] ), .B0(n2767), .Y(n2769) );
  AO21X1 U2531 ( .A0(n2766), .A1(n2765), .B0(n2764), .Y(n2767) );
  OAI21XL U2532 ( .A0(n2760), .A1(n2759), .B0(n2758), .Y(n2762) );
  OAI22XL U2533 ( .A0(n2755), .A1(n2754), .B0(n2757), .B1(\com[0][3] ), .Y(
        n2760) );
  INVX1 U2534 ( .A(n2261), .Y(n2262) );
  AOI211XL U2535 ( .A0(\com[1][1] ), .A1(n2752), .B0(n2751), .C0(\com[1][0] ), 
        .Y(n2755) );
  MXI2X2 U2536 ( .A(n2267), .B(n953), .S0(n1798), .Y(\com[1][1] ) );
  OAI22XL U2537 ( .A0(n2763), .A1(\com[0][4] ), .B0(\com[1][5] ), .B1(
        \com[0][5] ), .Y(n2765) );
  MXI2X2 U2538 ( .A(n2245), .B(n680), .S0(n1797), .Y(\com[0][7] ) );
  CLKINVX1 U2539 ( .A(n2251), .Y(n2253) );
  MXI2X2 U2540 ( .A(n2443), .B(n3240), .S0(n3126), .Y(n800) );
  MXI2X2 U2542 ( .A(n2442), .B(n3241), .S0(n3126), .Y(n795) );
  MXI2X2 U2546 ( .A(n2383), .B(n3244), .S0(n3126), .Y(n796) );
  NAND3X1 U2548 ( .A(n1800), .B(n3191), .C(n3190), .Y(n2440) );
  INVX1 U2550 ( .A(\com[3][0] ), .Y(n2365) );
  AO21X1 U2551 ( .A0(n2488), .A1(n2487), .B0(n2486), .Y(n2489) );
  NOR2X1 U2552 ( .A(\com[3][7] ), .B(n2485), .Y(n2364) );
  INVX1 U2553 ( .A(\com[2][2] ), .Y(n2353) );
  INVX1 U2554 ( .A(\com[2][0] ), .Y(n2351) );
  INVX1 U2555 ( .A(\com[2][1] ), .Y(n2352) );
  CLKINVX1 U2556 ( .A(n2582), .Y(n2349) );
  NAND2BX1 U2557 ( .AN(tree_mem_back[0]), .B(tree_mem_back[1]), .Y(n1818) );
  NAND2X1 U2558 ( .A(n2585), .B(n1720), .Y(n2330) );
  NAND3X4 U2560 ( .A(n2315), .B(n635), .C(\com[2][6] ), .Y(n2484) );
  INVX3 U2561 ( .A(n2314), .Y(n2315) );
  NAND3X2 U2562 ( .A(n2313), .B(n2487), .C(n2312), .Y(n2317) );
  NAND2X2 U2563 ( .A(n2477), .B(n2311), .Y(n2312) );
  NOR2X2 U2564 ( .A(\com[2][4] ), .B(n633), .Y(n2477) );
  NOR2X2 U2565 ( .A(n2310), .B(n2314), .Y(n2487) );
  NOR2X4 U2566 ( .A(\com[2][7] ), .B(n636), .Y(n2314) );
  OAI22X1 U2567 ( .A0(n635), .A1(\com[2][6] ), .B0(\com[2][5] ), .B1(n634), 
        .Y(n2310) );
  NAND2X2 U2568 ( .A(n2309), .B(n2480), .Y(n2313) );
  NAND2X1 U2569 ( .A(\com[2][4] ), .B(n633), .Y(n2308) );
  MXI2X4 U2570 ( .A(n2289), .B(n1761), .S0(n1780), .Y(\com[2][4] ) );
  NAND3X1 U2571 ( .A(n2306), .B(n2305), .C(n2478), .Y(n2482) );
  OAI21X1 U2572 ( .A0(n2476), .A1(n2479), .B0(n2478), .Y(n2307) );
  NAND2X1 U2573 ( .A(\com[2][3] ), .B(n632), .Y(n2478) );
  NOR2X1 U2574 ( .A(\com[2][2] ), .B(n631), .Y(n2479) );
  NOR2X1 U2575 ( .A(\com[2][3] ), .B(n632), .Y(n2476) );
  INVX3 U2576 ( .A(n2422), .Y(n2244) );
  NAND2X4 U2577 ( .A(\com[3][6] ), .B(n635), .Y(n2304) );
  CLKINVX1 U2578 ( .A(n2292), .Y(n2294) );
  MXI2X1 U2579 ( .A(n2620), .B(n2619), .S0(n1352), .Y(n2622) );
  NAND2X1 U2586 ( .A(state[2]), .B(n2946), .Y(n2951) );
  NOR2X1 U2587 ( .A(state[1]), .B(state[0]), .Y(n2946) );
  INVX3 U2590 ( .A(n2624), .Y(n2615) );
  INVX3 U2591 ( .A(n2447), .Y(n2599) );
  INVX4 U2592 ( .A(n2430), .Y(n2620) );
  NAND2X1 U2593 ( .A(n2426), .B(n2612), .Y(n2427) );
  OR2X4 U2594 ( .A(n2422), .B(n2421), .Y(n2430) );
  INVX3 U2595 ( .A(n2242), .Y(n2234) );
  NOR2X4 U2596 ( .A(n2418), .B(n2419), .Y(n2242) );
  INVX6 U2597 ( .A(n2421), .Y(n2402) );
  INVX3 U2598 ( .A(n1267), .Y(n2227) );
  MXI2X4 U2599 ( .A(n2415), .B(n2207), .S0(n1639), .Y(n2233) );
  INVX3 U2600 ( .A(n1304), .Y(n2207) );
  INVX3 U2601 ( .A(n1755), .Y(n2189) );
  INVX3 U2602 ( .A(n2263), .Y(n2178) );
  CLKINVX1 U2603 ( .A(n2270), .Y(n2170) );
  INVX1 U2604 ( .A(n2167), .Y(n2169) );
  CLKINVX1 U2605 ( .A(n949), .Y(n2166) );
  CLKINVX1 U2606 ( .A(n2293), .Y(n2202) );
  INVX3 U2607 ( .A(n2159), .Y(n2252) );
  MXI2X2 U2608 ( .A(n687), .B(n2250), .S0(n2152), .Y(n2268) );
  INVX3 U2609 ( .A(n2151), .Y(n2250) );
  INVX3 U2610 ( .A(n2259), .Y(n2182) );
  MXI2X4 U2611 ( .A(n680), .B(n2245), .S0(n2842), .Y(n2159) );
  INVX3 U2612 ( .A(n2130), .Y(n2245) );
  MXI2X4 U2613 ( .A(CNT6[4]), .B(n1391), .S0(n2152), .Y(n2259) );
  INVX3 U2614 ( .A(n2398), .Y(n2104) );
  INVX3 U2615 ( .A(n1301), .Y(n2095) );
  INVX1 U2616 ( .A(n2068), .Y(n2079) );
  INVX3 U2617 ( .A(n1997), .Y(n1994) );
  INVX3 U2618 ( .A(n1993), .Y(n1995) );
  INVX3 U2619 ( .A(n1990), .Y(n1991) );
  INVX3 U2620 ( .A(n2093), .Y(n1979) );
  INVX1 U2621 ( .A(n1337), .Y(n2083) );
  INVX4 U2622 ( .A(n2073), .Y(n2143) );
  INVX3 U2623 ( .A(n2040), .Y(n2115) );
  INVX3 U2624 ( .A(n2043), .Y(n2113) );
  MXI2X4 U2625 ( .A(n1944), .B(n1943), .S0(n1339), .Y(n2039) );
  INVX4 U2626 ( .A(n1981), .Y(n2058) );
  MXI2X4 U2627 ( .A(n1983), .B(n959), .S0(n1217), .Y(n1981) );
  INVX4 U2628 ( .A(n2057), .Y(n1982) );
  INVX3 U2629 ( .A(n1941), .Y(n1942) );
  INVX4 U2630 ( .A(n1943), .Y(n1946) );
  NOR2X4 U2631 ( .A(n1984), .B(n1950), .Y(n1941) );
  MXI2X4 U2632 ( .A(n1239), .B(n1230), .S0(n1325), .Y(n1944) );
  MXI2X4 U2633 ( .A(n1234), .B(n1171), .S0(n1325), .Y(n1950) );
  MXI2X4 U2634 ( .A(CNT3[6]), .B(n1930), .S0(n1025), .Y(n1984) );
  NAND2X6 U2635 ( .A(n2116), .B(CNT5[6]), .Y(n2031) );
  INVX6 U2636 ( .A(n2056), .Y(n2116) );
  MXI2X4 U2637 ( .A(n2014), .B(n673), .S0(n1786), .Y(n2056) );
  MXI2X4 U2638 ( .A(n1921), .B(n656), .S0(n1025), .Y(n1999) );
  CLKINVX1 U2639 ( .A(n659), .Y(n1926) );
  MXI2X4 U2640 ( .A(n1928), .B(CNT3[5]), .S0(n1137), .Y(n1915) );
  NAND2X6 U2641 ( .A(n1916), .B(CNT3[6]), .Y(n1909) );
  INVX6 U2642 ( .A(n1902), .Y(n1927) );
  MXI2X4 U2643 ( .A(n1171), .B(n1237), .S0(n1249), .Y(n1930) );
  NAND2X2 U2644 ( .A(n2585), .B(n3110), .Y(n2592) );
  OAI2BB1X1 U2645 ( .A0N(n2284), .A1N(N1142), .B0(n2276), .Y(n813) );
  INVX1 U2646 ( .A(\com[2][3] ), .Y(n2356) );
  INVX1 U2647 ( .A(n2415), .Y(n2416) );
  INVX2 U2648 ( .A(n1965), .Y(n2041) );
  MXI2X2 U2649 ( .A(n1211), .B(n1205), .S0(n1325), .Y(n1933) );
  INVX4 U2650 ( .A(n1910), .Y(n1921) );
  INVX1 U2651 ( .A(n1923), .Y(n1912) );
  INVX1 U2652 ( .A(\com[2][4] ), .Y(n2357) );
  INVX3 U2653 ( .A(n1947), .Y(n1948) );
  AOI21XL U2654 ( .A0(n2603), .A1(n611), .B0(n2602), .Y(n2604) );
  CLKINVX1 U2655 ( .A(n1324), .Y(n1898) );
  AOI211X1 U2656 ( .A0(n2479), .A1(n2478), .B0(n2477), .C0(n2476), .Y(n2481)
         );
  NAND2XL U2657 ( .A(n2700), .B(n1006), .Y(n2675) );
  MXI2XL U2658 ( .A(n2558), .B(n2557), .S0(n1012), .Y(n2659) );
  MXI2XL U2659 ( .A(n2571), .B(n2570), .S0(n1012), .Y(n2526) );
  MXI2X2 U2660 ( .A(n1250), .B(n2569), .S0(n998), .Y(n2684) );
  NAND2XL U2661 ( .A(n1798), .B(n1797), .Y(n2664) );
  MXI2XL U2662 ( .A(n2512), .B(n2511), .S0(n1796), .Y(n2574) );
  MXI2XL U2663 ( .A(n2497), .B(n2498), .S0(n972), .Y(n2506) );
  INVXL U2664 ( .A(n1326), .Y(n2493) );
  NAND2XL U2665 ( .A(n1006), .B(n2701), .Y(n2498) );
  MXI2XL U2666 ( .A(n2536), .B(n2537), .S0(n972), .Y(n2548) );
  MXI2XL U2667 ( .A(n2537), .B(n2536), .S0(n972), .Y(n2540) );
  AOI21XL U2668 ( .A0(n2531), .A1(n1326), .B0(n2530), .Y(n2536) );
  MXI2XL U2669 ( .A(n2571), .B(n2570), .S0(n1012), .Y(n2572) );
  INVXL U2670 ( .A(n1356), .Y(n2513) );
  INVX1 U2671 ( .A(n2925), .Y(n2923) );
  OAI21XL U2672 ( .A0(n2644), .A1(n775), .B0(n2643), .Y(n693) );
  INVX1 U2673 ( .A(n2913), .Y(n2934) );
  INVX1 U2674 ( .A(n2911), .Y(n2930) );
  OAI21XL U2675 ( .A0(tree_mem_back[1]), .A1(n1735), .B0(n2939), .Y(n2941) );
  OAI22XL U2676 ( .A0(n2935), .A1(n782), .B0(n2936), .B1(n1739), .Y(n777) );
  OAI21XL U2677 ( .A0(n1875), .A1(n680), .B0(n1874), .Y(n866) );
  NAND2X1 U2678 ( .A(n2911), .B(n1726), .Y(n2942) );
  OR3X1 U2679 ( .A(n1727), .B(tree_mem_back[1]), .C(tree_mem_back[0]), .Y(
        n1728) );
  NAND2X1 U2680 ( .A(n2757), .B(\com[0][3] ), .Y(n2758) );
  INVX1 U2681 ( .A(\com[1][3] ), .Y(n2757) );
  MXI2X2 U2682 ( .A(n2263), .B(n2262), .S0(n1798), .Y(\com[1][3] ) );
  MXI2X4 U2683 ( .A(n2270), .B(n2269), .S0(n1798), .Y(\com[1][0] ) );
  INVX1 U2685 ( .A(n2448), .Y(n2438) );
  NAND2BXL U2686 ( .AN(n3109), .B(n3110), .Y(n2321) );
  INVX1 U2687 ( .A(n1781), .Y(n2332) );
  OAI2BB1X1 U2691 ( .A0N(n802), .A1N(n636), .B0(n2348), .Y(n2582) );
  NAND2X1 U2692 ( .A(n2913), .B(n810), .Y(n2933) );
  NAND2XL U2693 ( .A(tree_mem_back[1]), .B(tree_mem_back[0]), .Y(n1817) );
  MXI2X4 U2694 ( .A(n1296), .B(n977), .S0(n930), .Y(n2596) );
  MXI2X4 U2695 ( .A(n2412), .B(n2411), .S0(n1796), .Y(n2435) );
  MXI2X4 U2696 ( .A(n2408), .B(n2407), .S0(n1796), .Y(n2597) );
  MXI2X4 U2697 ( .A(n2393), .B(n975), .S0(n1801), .Y(n2601) );
  MXI2X4 U2698 ( .A(n1567), .B(n1314), .S0(n1639), .Y(n2275) );
  MXI2X4 U2699 ( .A(n1762), .B(n1014), .S0(n1494), .Y(n2208) );
  MXI2X4 U2700 ( .A(n2261), .B(n2178), .S0(n1474), .Y(n2295) );
  MXI2X4 U2701 ( .A(n2140), .B(n2139), .S0(n1791), .Y(n2181) );
  MXI2X4 U2702 ( .A(n2391), .B(n2390), .S0(n1796), .Y(n2600) );
  AND2X8 U2703 ( .A(n2108), .B(n2107), .Y(n2398) );
  MXI2X4 U2704 ( .A(n2095), .B(n1755), .S0(n1793), .Y(n2225) );
  MXI2X2 U2705 ( .A(n2080), .B(n2079), .S0(n1788), .Y(n2203) );
  MXI2X4 U2706 ( .A(n1168), .B(n2093), .S0(n1788), .Y(n2213) );
  MXI2X4 U2707 ( .A(n1774), .B(n2086), .S0(n1788), .Y(n2411) );
  MXI2X4 U2708 ( .A(n676), .B(n964), .S0(n1786), .Y(n2046) );
  INVX3 U2709 ( .A(n1934), .Y(n1977) );
  MXI2X4 U2710 ( .A(CNT3[3]), .B(n1927), .S0(n1137), .Y(n1935) );
  MXI2X4 U2711 ( .A(n2001), .B(CNT4[5]), .S0(n1786), .Y(n2013) );
  MXI2X4 U2712 ( .A(n1064), .B(n678), .S0(n1786), .Y(n2051) );
  MXI2X4 U2713 ( .A(n1204), .B(n1210), .S0(n1249), .Y(n1911) );
  OAI21X4 U2714 ( .A0(n1890), .A1(n1891), .B0(n1889), .Y(n1897) );
  OAI21X4 U2715 ( .A0(n1888), .A1(n1887), .B0(n1886), .Y(n1889) );
  OAI21X4 U2716 ( .A0(n1882), .A1(n1883), .B0(n1881), .Y(n1891) );
  NAND2BX4 U2717 ( .AN(n1210), .B(n1204), .Y(n1880) );
  CLKBUFX3 U2719 ( .A(n1805), .Y(n1807) );
  CLKBUFX3 U2720 ( .A(n1806), .Y(n1805) );
  CLKBUFX3 U2721 ( .A(n2914), .Y(n1806) );
  CLKBUFX3 U2725 ( .A(n1804), .Y(n1811) );
  CLKBUFX3 U2726 ( .A(n2914), .Y(n1804) );
  AND4X1 U2728 ( .A(n2785), .B(n2957), .C(n2784), .D(n2783), .Y(n2786) );
  AOI22X1 U2729 ( .A0(n1134), .A1(n3059), .B0(n2743), .B1(n3060), .Y(n3036) );
  OAI22XL U2730 ( .A0(n2852), .A1(n1115), .B0(n2851), .B1(n1703), .Y(N682) );
  OAI22XL U2731 ( .A0(n2860), .A1(n1115), .B0(n1703), .B1(n2859), .Y(N724) );
  AOI22XL U2732 ( .A0(n3053), .A1(n2843), .B0(n3052), .B1(n1797), .Y(n2845) );
  AOI22XL U2733 ( .A0(n3056), .A1(n2843), .B0(n3055), .B1(n1797), .Y(n2841) );
  OAI21XL U2734 ( .A0(n1723), .A1(n2952), .B0(n2953), .Y(N720) );
  OAI22XL U2735 ( .A0(n2850), .A1(n1115), .B0(n2849), .B1(n1703), .Y(N668) );
  OAI22XL U2736 ( .A0(n2856), .A1(n1115), .B0(n2855), .B1(n1703), .Y(N710) );
  OAI22XL U2737 ( .A0(n2848), .A1(n1703), .B0(n2847), .B1(n1115), .Y(N654) );
  OAI22XL U2738 ( .A0(n2854), .A1(n1115), .B0(n2853), .B1(n1703), .Y(N696) );
  OAI222XL U2739 ( .A0(n1694), .A1(n2829), .B0(n1097), .B1(n2854), .C0(n2853), 
        .C1(n1114), .Y(N690) );
  OAI22XL U2740 ( .A0(n2854), .A1(n1096), .B0(n2853), .B1(n1113), .Y(N691) );
  OR2X2 U2741 ( .A(n2709), .B(n2715), .Y(n2853) );
  AOI22XL U2742 ( .A0(n3067), .A1(n2843), .B0(n3066), .B1(n1797), .Y(n2832) );
  OAI222XL U2743 ( .A0(n1694), .A1(n2828), .B0(n1097), .B1(n2852), .C0(n2851), 
        .C1(n1114), .Y(N676) );
  INVX1 U2744 ( .A(n3020), .Y(n2713) );
  OAI222XL U2745 ( .A0(n1114), .A1(n2859), .B0(n1097), .B1(n2860), .C0(n1694), 
        .C1(n2858), .Y(N718) );
  AOI22X1 U2746 ( .A0(n1134), .A1(n3070), .B0(n2743), .B1(n3071), .Y(n3043) );
  INVX1 U2747 ( .A(n2705), .Y(n2788) );
  INVX1 U2748 ( .A(n3040), .Y(n2775) );
  OAI222XL U2749 ( .A0(n1694), .A1(n2830), .B0(n1097), .B1(n2856), .C0(n2855), 
        .C1(n1114), .Y(N704) );
  OAI22XL U2750 ( .A0(n2848), .A1(n1113), .B0(n2847), .B1(n1096), .Y(N649) );
  INVX1 U2751 ( .A(n1134), .Y(n2848) );
  OAI211X1 U2752 ( .A0(n2721), .A1(n3020), .B0(n3045), .C0(n2960), .Y(n2704)
         );
  INVX1 U2753 ( .A(n2959), .Y(n2724) );
  NAND2BX1 U2754 ( .AN(n3018), .B(n2796), .Y(n3002) );
  INVX1 U2755 ( .A(n2721), .Y(n2714) );
  OAI21XL U2756 ( .A0(n2909), .A1(n3019), .B0(n2900), .Y(n3018) );
  OAI22XL U2757 ( .A0(n2852), .A1(n1096), .B0(n2851), .B1(n1113), .Y(N677) );
  INVX1 U2758 ( .A(n2901), .Y(n2851) );
  OAI222XL U2759 ( .A0(n1114), .A1(n2849), .B0(n1097), .B1(n2850), .C0(n2827), 
        .C1(n1694), .Y(N662) );
  OR2X2 U2760 ( .A(n1797), .B(n2702), .Y(n2847) );
  OR2X2 U2761 ( .A(n1797), .B(n2696), .Y(n2852) );
  NOR2XL U2762 ( .A(n1797), .B(n1323), .Y(n2700) );
  OR2X2 U2763 ( .A(n1797), .B(n2679), .Y(n2854) );
  OAI22XL U2764 ( .A0(n2856), .A1(n1096), .B0(n2855), .B1(n1113), .Y(N705) );
  OR2X2 U2765 ( .A(n1797), .B(n2668), .Y(n2856) );
  OAI22XL U2766 ( .A0(n2860), .A1(n1096), .B0(n1113), .B1(n2859), .Y(N719) );
  OAI22XL U2767 ( .A0(n2850), .A1(n1096), .B0(n2849), .B1(n1113), .Y(N663) );
  OAI2BB1X1 U2768 ( .A0N(n1265), .A1N(n2667), .B0(n2666), .Y(n2715) );
  MXI2XL U2769 ( .A(n2545), .B(n2544), .S0(n1796), .Y(n2660) );
  OR2X1 U2770 ( .A(n2960), .B(n2655), .Y(n2846) );
  AND2X1 U2771 ( .A(n2859), .B(n2860), .Y(n2652) );
  INVX1 U2772 ( .A(n2703), .Y(n2718) );
  INVX1 U2773 ( .A(n2565), .Y(n2568) );
  INVX1 U2774 ( .A(n2561), .Y(n2564) );
  AND2X1 U2775 ( .A(n2960), .B(n1743), .Y(n2998) );
  OAI22XL U2776 ( .A0(n2508), .A1(n2695), .B0(n1265), .B1(n2507), .Y(n2562) );
  NOR2X1 U2777 ( .A(n1058), .B(n2504), .Y(n2695) );
  AND2X1 U2778 ( .A(n2523), .B(n2496), .Y(n2510) );
  NOR2X1 U2779 ( .A(n1326), .B(n1325), .Y(n2504) );
  OR2X1 U2780 ( .A(n2720), .B(n2721), .Y(n2960) );
  OR2X1 U2781 ( .A(n1323), .B(n2546), .Y(n2694) );
  MXI2XL U2782 ( .A(n2553), .B(n2552), .S0(n1796), .Y(n2557) );
  AND2X1 U2783 ( .A(n1323), .B(n2527), .Y(n2547) );
  NOR2XL U2784 ( .A(n1006), .B(n2532), .Y(n2546) );
  NOR2XL U2785 ( .A(n1326), .B(n2534), .Y(n2532) );
  INVXL U2786 ( .A(n1325), .Y(n2534) );
  CLKINVX2 U2787 ( .A(n1797), .Y(n2860) );
  XOR2XL U2788 ( .A(n2322), .B(n3109), .Y(n1815) );
  OAI21XL U2789 ( .A0(n2938), .A1(n2865), .B0(n2641), .Y(n696) );
  OAI21XL U2790 ( .A0(n2585), .A1(n1720), .B0(n1781), .Y(n820) );
  OAI22XL U2791 ( .A0(n2642), .A1(n775), .B0(n2913), .B1(n1714), .Y(n774) );
  OAI21XL U2792 ( .A0(n1714), .A1(n2935), .B0(n2584), .Y(n773) );
  OAI21XL U2793 ( .A0(n579), .A1(n2943), .B0(n2944), .Y(n755) );
  OAI21XL U2794 ( .A0(n1783), .A1(n1214), .B0(n1843), .Y(n841) );
  OAI21XL U2795 ( .A0(n1783), .A1(n1239), .B0(n1844), .Y(n834) );
  OAI21XL U2796 ( .A0(n1783), .A1(n1211), .B0(n1839), .Y(n837) );
  OAI21XL U2797 ( .A0(n1783), .A1(n1199), .B0(n1840), .Y(n838) );
  OAI21XL U2798 ( .A0(n1783), .A1(n1475), .B0(n1842), .Y(n840) );
  OAI21XL U2799 ( .A0(n1783), .A1(n1208), .B0(n1838), .Y(n836) );
  OAI21XL U2800 ( .A0(n1783), .A1(n1237), .B0(n1837), .Y(n835) );
  OAI21XL U2801 ( .A0(n1783), .A1(n1885), .B0(n1841), .Y(n839) );
  OAI21XL U2802 ( .A0(n1782), .A1(n679), .B0(n1825), .Y(n865) );
  OAI21XL U2803 ( .A0(n1782), .A1(n672), .B0(n1826), .Y(n858) );
  OAI21XL U2804 ( .A0(n1782), .A1(n677), .B0(n1823), .Y(n863) );
  OAI21XL U2805 ( .A0(n1782), .A1(n673), .B0(n1819), .Y(n859) );
  OAI21XL U2806 ( .A0(n1782), .A1(n675), .B0(n1821), .Y(n861) );
  OAI21XL U2807 ( .A0(n1782), .A1(n674), .B0(n1820), .Y(n860) );
  OAI21XL U2808 ( .A0(n1782), .A1(n676), .B0(n1822), .Y(n862) );
  OAI21XL U2809 ( .A0(n1782), .A1(n678), .B0(n1824), .Y(n864) );
  MXI2X2 U2810 ( .A(n2247), .B(n683), .S0(n1797), .Y(\com[0][4] ) );
  OAI2BB1X4 U2811 ( .A0N(n2304), .A1N(n2316), .B0(\com[3][7] ), .Y(n2320) );
  MXI2X4 U2812 ( .A(n2294), .B(n2293), .S0(n1780), .Y(\com[2][1] ) );
  OR2X2 U2813 ( .A(n2929), .B(n1816), .Y(n2938) );
  NAND2BXL U2814 ( .AN(tree_mem_back[1]), .B(tree_mem_back[0]), .Y(n1816) );
  MXI2X4 U2815 ( .A(n2619), .B(n2620), .S0(n1352), .Y(\com[4][7] ) );
  MXI2X4 U2816 ( .A(n2599), .B(n2601), .S0(n1803), .Y(\com[4][0] ) );
  MXI2X4 U2817 ( .A(n1481), .B(n2132), .S0(n1648), .Y(n2251) );
  MXI2X4 U2818 ( .A(n2109), .B(n664), .S0(n1323), .Y(n2130) );
  MXI2X4 U2819 ( .A(CNT4[6]), .B(n1949), .S0(n1279), .Y(n2057) );
  MXI2X2 U2820 ( .A(n1208), .B(n1766), .S0(n1325), .Y(n1931) );
  MXI2X2 U2821 ( .A(n1199), .B(n1324), .S0(n1343), .Y(n1971) );
  MXI2X4 U2822 ( .A(n1590), .B(n672), .S0(n1336), .Y(n2034) );
  NAND2BX4 U2823 ( .AN(n1229), .B(n1238), .Y(n1892) );
  NOR3X1 U2825 ( .A(n2782), .B(n2781), .C(n2780), .Y(n2785) );
  INVX1 U2826 ( .A(n2849), .Y(n2780) );
  NOR3X1 U2827 ( .A(n2903), .B(n2689), .C(n2688), .Y(n2690) );
  INVX1 U2828 ( .A(n2853), .Y(n2688) );
  INVX1 U2829 ( .A(n2854), .Y(n2689) );
  AOI211X1 U2830 ( .A0(n2986), .A1(n3000), .B0(n2902), .C0(n3001), .Y(n2999)
         );
  INVX1 U2831 ( .A(n2985), .Y(n3001) );
  INVX1 U2832 ( .A(n2691), .Y(n2692) );
  OAI211X1 U2833 ( .A0(n2746), .A1(n2745), .B0(n2799), .C0(n2744), .Y(n2748)
         );
  INVX1 U2834 ( .A(n2904), .Y(n2744) );
  AOI211X1 U2835 ( .A0(n2982), .A1(n2983), .B0(n2905), .C0(n2979), .Y(n2978)
         );
  OAI211X1 U2836 ( .A0(n2984), .A1(n2957), .B0(n2985), .C0(n2977), .Y(n2983)
         );
  NOR2X1 U2837 ( .A(n2998), .B(n2955), .Y(n2985) );
  AOI211X1 U2838 ( .A0(n2579), .A1(n2693), .B0(n2998), .C0(n2578), .Y(n2580)
         );
  NAND4X1 U2839 ( .A(n2860), .B(n2956), .C(n2954), .D(n2859), .Y(n2578) );
  INVX1 U2840 ( .A(n2960), .Y(n2579) );
  INVX1 U2841 ( .A(n2955), .Y(n2581) );
  INVX1 U2842 ( .A(n2804), .Y(n2554) );
  OR4X2 U2843 ( .A(n2806), .B(n2805), .C(n2804), .D(n2803), .Y(N672) );
  OAI211X1 U2844 ( .A0(n2802), .A1(n2801), .B0(n2800), .C0(n2799), .Y(n2803)
         );
  INVX1 U2845 ( .A(n2998), .Y(n2799) );
  AOI211X1 U2846 ( .A0(n2798), .A1(n2797), .B0(n2796), .C0(n2795), .Y(n2800)
         );
  NAND2X1 U2847 ( .A(n2852), .B(n2851), .Y(n2795) );
  NOR2X1 U2848 ( .A(n2745), .B(n2783), .Y(n2804) );
  NAND2X1 U2849 ( .A(n2736), .B(n2801), .Y(n2783) );
  INVX1 U2850 ( .A(n2957), .Y(n2806) );
  OAI211X1 U2851 ( .A0(n2705), .A1(n2684), .B0(n2685), .C0(n2787), .Y(n2957)
         );
  NAND2X1 U2852 ( .A(n3047), .B(n3048), .Y(N203) );
  NAND2X1 U2853 ( .A(n2743), .B(n3052), .Y(n3033) );
  NAND2X1 U2854 ( .A(n2743), .B(n3055), .Y(n3035) );
  AOI31X1 U2855 ( .A0(n2777), .A1(n2776), .A2(n3061), .B0(n2742), .Y(n3039) );
  OAI211X1 U2856 ( .A0(n1731), .A1(n3038), .B0(n2741), .C0(n2740), .Y(n2742)
         );
  AOI2BB2X1 U2857 ( .B0(n2743), .B1(n3063), .A0N(n1693), .A1N(n2848), .Y(n2741) );
  NAND2X1 U2858 ( .A(n2899), .B(n3051), .Y(n3004) );
  AOI2BB2X1 U2859 ( .B0(n2901), .B1(n3053), .A0N(n2852), .A1N(n1697), .Y(n3003) );
  NAND2X1 U2860 ( .A(n2899), .B(n3054), .Y(n3006) );
  AOI2BB2X1 U2861 ( .B0(n2901), .B1(n3056), .A0N(n2852), .A1N(n1698), .Y(n3005) );
  AOI2BB2X1 U2862 ( .B0(n2899), .B1(n3058), .A0N(n3009), .A1N(n1713), .Y(n3008) );
  AOI2BB2X1 U2863 ( .B0(n2901), .B1(n3059), .A0N(n2852), .A1N(n1118), .Y(n3007) );
  AOI211X1 U2864 ( .A0(n2901), .A1(n3050), .B0(n3011), .C0(n3012), .Y(n3010)
         );
  NAND2X1 U2865 ( .A(n2837), .B(n3057), .Y(n2838) );
  AOI211X1 U2866 ( .A0(n2857), .A1(n3062), .B0(n2657), .C0(n2656), .Y(n2658)
         );
  NOR2X1 U2867 ( .A(n1730), .B(n2846), .Y(n2657) );
  NAND2X1 U2868 ( .A(n2898), .B(n3051), .Y(n3022) );
  NAND2X1 U2869 ( .A(n2898), .B(n3054), .Y(n3023) );
  AOI2BB2X1 U2870 ( .B0(n2898), .B1(n3058), .A0N(n3025), .A1N(n1713), .Y(n3024) );
  OA22X1 U2871 ( .A0(n2849), .A1(n1705), .B0(n2850), .B1(n1118), .Y(n1746) );
  AOI211X1 U2872 ( .A0(n3063), .A1(n2782), .B0(n2725), .C0(n3027), .Y(n2726)
         );
  NOR2X1 U2873 ( .A(n1693), .B(n2849), .Y(n2725) );
  NAND2X1 U2874 ( .A(n2905), .B(n3051), .Y(n2963) );
  OA22X1 U2875 ( .A0(n2856), .A1(n1697), .B0(n2855), .B1(n1708), .Y(n2962) );
  NAND2X1 U2876 ( .A(n2905), .B(n3054), .Y(n2965) );
  OA22X1 U2877 ( .A0(n2856), .A1(n1698), .B0(n2855), .B1(n1709), .Y(n2964) );
  AOI211X1 U2878 ( .A0(n2905), .A1(n3062), .B0(n2970), .C0(n2971), .Y(n2969)
         );
  NAND2X1 U2879 ( .A(n2903), .B(n3051), .Y(n2988) );
  NAND2X1 U2880 ( .A(n2903), .B(n3054), .Y(n2989) );
  AOI2BB2X1 U2881 ( .B0(n2903), .B1(n3058), .A0N(n2991), .A1N(n1713), .Y(n2990) );
  AOI211X1 U2882 ( .A0(n3062), .A1(n2903), .B0(n2993), .C0(n2994), .Y(n2992)
         );
  AOI2BB2X1 U2883 ( .B0(n2903), .B1(n3069), .A0N(n2991), .A1N(n1733), .Y(n2997) );
  NAND2X1 U2884 ( .A(n2903), .B(n3064), .Y(n2996) );
  INVX1 U2885 ( .A(n2903), .Y(n2829) );
  OAI211X1 U2886 ( .A0(n2995), .A1(n1742), .B0(n2816), .C0(n2815), .Y(N687) );
  NAND2X1 U2887 ( .A(n775), .B(n2814), .Y(n2815) );
  INVX1 U2888 ( .A(n2991), .Y(n2814) );
  NAND3X1 U2889 ( .A(n2802), .B(n2691), .C(n2687), .Y(n2991) );
  INVX1 U2890 ( .A(n2745), .Y(n2802) );
  AOI211X1 U2891 ( .A0(n776), .A1(n2903), .B0(n2813), .C0(n2812), .Y(n2816) );
  NAND2X1 U2892 ( .A(n2683), .B(n2676), .Y(n2677) );
  INVX1 U2893 ( .A(n2682), .Y(n2676) );
  NOR2X2 U2894 ( .A(n2681), .B(n2680), .Y(n2903) );
  NAND2X1 U2895 ( .A(n2687), .B(n2902), .Y(n2995) );
  AOI211X1 U2896 ( .A0(n2686), .A1(n2958), .B0(n2685), .C0(n2684), .Y(n2902)
         );
  NAND2X1 U2897 ( .A(n2705), .B(n2671), .Y(n2685) );
  NOR2X1 U2898 ( .A(n2724), .B(n2734), .Y(n2686) );
  AOI211X1 U2899 ( .A0(n2714), .A1(n2683), .B0(n2998), .C0(n2682), .Y(n2687)
         );
  NAND2X1 U2900 ( .A(n2853), .B(n2675), .Y(n2680) );
  NAND2X1 U2901 ( .A(n2837), .B(n3068), .Y(n2834) );
  OAI211X1 U2902 ( .A0(n2966), .A1(n1733), .B0(n2975), .C0(n2976), .Y(N702) );
  OA22X1 U2903 ( .A0(n1706), .A1(n2855), .B0(n1696), .B1(n2856), .Y(n2975) );
  NAND2X1 U2904 ( .A(n2857), .B(n3064), .Y(n2831) );
  INVX1 U2905 ( .A(n2859), .Y(n2843) );
  OA22X1 U2906 ( .A0(n2856), .A1(n1707), .B0(n2855), .B1(n1699), .Y(n2973) );
  OAI211X1 U2907 ( .A0(n2966), .A1(n1713), .B0(n2967), .C0(n2968), .Y(N707) );
  OA22X1 U2908 ( .A0(n1705), .A1(n2855), .B0(n1118), .B1(n2856), .Y(n2967) );
  OAI211X1 U2909 ( .A0(n2972), .A1(n1742), .B0(n2821), .C0(n2820), .Y(N701) );
  NAND2X1 U2910 ( .A(n775), .B(n2819), .Y(n2820) );
  INVX1 U2911 ( .A(n2966), .Y(n2819) );
  NAND3X1 U2912 ( .A(n2734), .B(n2672), .C(n2746), .Y(n2966) );
  INVX1 U2913 ( .A(n2736), .Y(n2746) );
  INVX1 U2915 ( .A(n2979), .Y(n2669) );
  NAND2BX1 U2916 ( .AN(n2977), .B(n2672), .Y(n2972) );
  NOR2X1 U2917 ( .A(n2979), .B(n2980), .Y(n2672) );
  NAND2X1 U2918 ( .A(n2907), .B(n2954), .Y(n2982) );
  INVX1 U2919 ( .A(n2674), .Y(n2907) );
  NAND3BX1 U2920 ( .AN(n2984), .B(n2671), .C(n2788), .Y(n2977) );
  NAND2X1 U2921 ( .A(n2906), .B(n2959), .Y(n2986) );
  INVX1 U2922 ( .A(n2899), .Y(n2828) );
  NAND2X1 U2923 ( .A(n2899), .B(n3064), .Y(n3015) );
  AOI2BB2X1 U2924 ( .B0(n2901), .B1(n3067), .A0N(n2852), .A1N(n1707), .Y(n3014) );
  NAND2X1 U2925 ( .A(n2898), .B(n3064), .Y(n3029) );
  OAI211X1 U2926 ( .A0(n3028), .A1(n1742), .B0(n2794), .C0(n2793), .Y(N659) );
  NAND2X1 U2927 ( .A(n775), .B(n2792), .Y(n2793) );
  INVX1 U2928 ( .A(n3025), .Y(n2792) );
  NAND3BX1 U2929 ( .AN(n2727), .B(n2724), .C(n2801), .Y(n3025) );
  AOI211X1 U2930 ( .A0(n776), .A1(n2898), .B0(n2791), .C0(n2790), .Y(n2794) );
  NAND3X1 U2931 ( .A(n2714), .B(n2713), .C(n2722), .Y(n3021) );
  OR4X1 U2932 ( .A(n2789), .B(n2787), .C(n2788), .D(n2727), .Y(n3028) );
  NAND3X1 U2933 ( .A(n2723), .B(n2722), .C(n2784), .Y(n2727) );
  NAND2BX1 U2934 ( .AN(n2721), .B(n2720), .Y(n2784) );
  NOR2X1 U2935 ( .A(n2781), .B(n2717), .Y(n2722) );
  NOR2X1 U2936 ( .A(n2798), .B(n2732), .Y(n2781) );
  NAND2X1 U2937 ( .A(n2719), .B(n2721), .Y(n2723) );
  OAI211X1 U2938 ( .A0(n3013), .A1(n1742), .B0(n2811), .C0(n2810), .Y(N673) );
  NAND2X1 U2939 ( .A(n775), .B(n2809), .Y(n2810) );
  INVX1 U2940 ( .A(n3009), .Y(n2809) );
  AOI211X1 U2941 ( .A0(n776), .A1(n2899), .B0(n2808), .C0(n2807), .Y(n2811) );
  NAND2X1 U2942 ( .A(n2707), .B(n2805), .Y(n3013) );
  AOI211X1 U2943 ( .A0(n2906), .A1(n2706), .B0(n2705), .C0(n2787), .Y(n2805)
         );
  NAND2X1 U2944 ( .A(n2737), .B(n2684), .Y(n2787) );
  NAND2X1 U2945 ( .A(n2724), .B(n2801), .Y(n2706) );
  OAI211X1 U2946 ( .A0(n3031), .A1(n1717), .B0(n3041), .C0(n3042), .Y(N647) );
  NAND2X1 U2947 ( .A(n2743), .B(n3066), .Y(n3042) );
  INVX1 U2948 ( .A(n2857), .Y(n2858) );
  INVX1 U2949 ( .A(n2847), .Y(n2743) );
  OAI211X1 U2950 ( .A0(n1719), .A1(n3038), .B0(n2779), .C0(n2778), .Y(N645) );
  NAND3X1 U2951 ( .A(n2777), .B(n2865), .C(n2776), .Y(n2778) );
  MXI2X1 U2952 ( .A(n2663), .B(n2662), .S0(n998), .Y(n2705) );
  INVX1 U2953 ( .A(n2660), .Y(n2662) );
  INVX1 U2954 ( .A(n2659), .Y(n2663) );
  NOR2X1 U2955 ( .A(n2691), .B(n2734), .Y(n2906) );
  INVX1 U2956 ( .A(n2684), .Y(n2739) );
  AOI211X1 U2957 ( .A0(n776), .A1(n2775), .B0(n2774), .C0(n2773), .Y(n2779) );
  NAND2X1 U2958 ( .A(n2747), .B(n2904), .Y(n3031) );
  NOR2X1 U2959 ( .A(n2673), .B(n3045), .Y(n2904) );
  INVX1 U2960 ( .A(n2720), .Y(n2673) );
  NAND3X1 U2961 ( .A(n2736), .B(n2734), .C(n2776), .Y(n3038) );
  AOI2BB1X1 U2962 ( .A0N(n2732), .A1N(n2797), .B0(n2731), .Y(n2747) );
  INVX1 U2963 ( .A(n2735), .Y(n2731) );
  INVX1 U2964 ( .A(n2728), .Y(n2797) );
  NAND2X1 U2965 ( .A(n2960), .B(n3020), .Y(n2981) );
  NOR2X1 U2966 ( .A(n2720), .B(n3045), .Y(n2733) );
  NOR2X1 U2967 ( .A(n2801), .B(n2745), .Y(n2734) );
  NAND2X1 U2968 ( .A(n2735), .B(n2909), .Y(n3040) );
  AOI2BB2X1 U2969 ( .B0(n2730), .B1(n2852), .A0N(n2901), .A1N(n2729), .Y(n2735) );
  INVX1 U2970 ( .A(n2905), .Y(n2830) );
  NOR3X2 U2971 ( .A(n2708), .B(n2670), .C(n2979), .Y(n2905) );
  NAND2X1 U2972 ( .A(n2855), .B(n2856), .Y(n2979) );
  NAND3X1 U2973 ( .A(n2724), .B(n2707), .C(n1251), .Y(n3009) );
  NOR2BX1 U2974 ( .AN(n2704), .B(n3018), .Y(n2707) );
  NAND2X1 U2975 ( .A(n2736), .B(n2745), .Y(n2959) );
  AND3X2 U2976 ( .A(n2798), .B(n2703), .C(n2900), .Y(n2899) );
  AOI2BB2X1 U2977 ( .B0(n2901), .B1(n3070), .A0N(n2852), .A1N(n1696), .Y(n3016) );
  NOR2X1 U2978 ( .A(n2714), .B(n3020), .Y(n2796) );
  AOI2BB2X1 U2979 ( .B0(n2730), .B1(n2847), .A0N(n1134), .A1N(n2729), .Y(n2900) );
  NAND2X1 U2980 ( .A(n2715), .B(n2710), .Y(n2729) );
  NOR2X1 U2981 ( .A(n2782), .B(n2712), .Y(n2730) );
  MXI2X1 U2982 ( .A(n2798), .B(n2708), .S0(n2728), .Y(n3019) );
  INVX1 U2983 ( .A(n2732), .Y(n2708) );
  INVX1 U2984 ( .A(n2898), .Y(n2827) );
  NOR3X2 U2985 ( .A(n2798), .B(n2718), .C(n2717), .Y(n2898) );
  NAND2X1 U2986 ( .A(n2852), .B(n2847), .Y(n2711) );
  NAND2X1 U2987 ( .A(n2695), .B(n2694), .Y(n2696) );
  NAND2X1 U2988 ( .A(n2854), .B(n2700), .Y(n2712) );
  NAND2X1 U2989 ( .A(n2678), .B(n2697), .Y(n2679) );
  INVX1 U2990 ( .A(n2695), .Y(n2678) );
  AND2X2 U2991 ( .A(n2709), .B(n2715), .Y(n2901) );
  NAND2BX2 U2992 ( .AN(n2710), .B(n2715), .Y(n2855) );
  OR2X2 U2993 ( .A(n2716), .B(n2715), .Y(n2849) );
  NAND2X1 U2994 ( .A(n2665), .B(n2694), .Y(n2666) );
  INVX1 U2995 ( .A(n2664), .Y(n2665) );
  NAND2X1 U2996 ( .A(n2710), .B(n2709), .Y(n2716) );
  NOR2X1 U2997 ( .A(n1797), .B(n2699), .Y(n2782) );
  NAND2X1 U2998 ( .A(n2698), .B(n2697), .Y(n2699) );
  INVX1 U2999 ( .A(n2694), .Y(n2697) );
  OAI211X1 U3000 ( .A0(n1742), .A1(n2952), .B0(n2826), .C0(n2825), .Y(N715) );
  NAND2X1 U3001 ( .A(n775), .B(n2837), .Y(n2825) );
  INVX1 U3002 ( .A(n2824), .Y(n2837) );
  NAND2X1 U3003 ( .A(n2651), .B(n2650), .Y(n2824) );
  INVX1 U3004 ( .A(n2958), .Y(n2651) );
  NAND2X1 U3005 ( .A(n2691), .B(n2745), .Y(n2958) );
  MXI2X2 U3006 ( .A(n2569), .B(n1250), .S0(n998), .Y(n2745) );
  NOR2X1 U3007 ( .A(n2736), .B(n1251), .Y(n2691) );
  INVX1 U3008 ( .A(n2553), .Y(n2544) );
  MXI2X1 U3009 ( .A(n2539), .B(n2538), .S0(n1794), .Y(n2545) );
  INVX1 U3010 ( .A(n2646), .Y(n2538) );
  INVX1 U3011 ( .A(n2645), .Y(n2539) );
  MXI2X2 U3012 ( .A(n1120), .B(n2526), .S0(n998), .Y(n2736) );
  AOI211X1 U3013 ( .A0(n776), .A1(n2857), .B0(n2823), .C0(n2822), .Y(n2826) );
  INVX1 U3014 ( .A(n2652), .Y(n2653) );
  NAND2BX1 U3015 ( .AN(n2728), .B(n2732), .Y(n2954) );
  NAND3X1 U3016 ( .A(n2671), .B(n2650), .C(n2684), .Y(n2952) );
  INVX1 U3017 ( .A(n2512), .Y(n2502) );
  INVX1 U3018 ( .A(n2511), .Y(n2503) );
  NOR3X1 U3019 ( .A(n2998), .B(n2719), .C(n2654), .Y(n2650) );
  NAND2BX2 U3020 ( .AN(n2710), .B(n2709), .Y(n2859) );
  OAI22X1 U3021 ( .A0(n2664), .A1(n1058), .B0(n1798), .B1(n2575), .Y(n2710) );
  INVX1 U3022 ( .A(n2670), .Y(n2649) );
  NAND3X1 U3023 ( .A(n2648), .B(n2718), .C(n2681), .Y(n2674) );
  NAND2X1 U3024 ( .A(n2908), .B(n2732), .Y(n2681) );
  NOR2BX1 U3025 ( .AN(n2728), .B(n2798), .Y(n2908) );
  NOR2X1 U3026 ( .A(n2728), .B(n2732), .Y(n2703) );
  INVX1 U3027 ( .A(n2909), .Y(n2648) );
  NOR2X1 U3028 ( .A(n2670), .B(n2732), .Y(n2909) );
  MXI2X2 U3029 ( .A(n2568), .B(n2567), .S0(n1780), .Y(n2732) );
  INVX1 U3030 ( .A(n2566), .Y(n2567) );
  NAND2X1 U3031 ( .A(n2728), .B(n2798), .Y(n2670) );
  MXI2X2 U3032 ( .A(n2551), .B(n2647), .S0(n1780), .Y(n2798) );
  MXI2X2 U3033 ( .A(n2564), .B(n2563), .S0(n1780), .Y(n2728) );
  INVX1 U3034 ( .A(n2562), .Y(n2563) );
  NOR2X1 U3035 ( .A(n2720), .B(n2683), .Y(n2719) );
  NAND2X1 U3036 ( .A(n2720), .B(n2693), .Y(n3020) );
  INVX1 U3037 ( .A(n2683), .Y(n2693) );
  NAND2X1 U3038 ( .A(n2683), .B(n2721), .Y(n3045) );
  MXI2X2 U3039 ( .A(n2574), .B(n2573), .S0(n995), .Y(n2683) );
  MXI2X1 U3040 ( .A(n2510), .B(n2509), .S0(n1794), .Y(n2561) );
  INVX1 U3041 ( .A(n2577), .Y(n2507) );
  MXI2X1 U3042 ( .A(n2506), .B(n2505), .S0(n1008), .Y(n2577) );
  INVX1 U3043 ( .A(n2550), .Y(n2508) );
  MXI2X1 U3044 ( .A(n2509), .B(n2510), .S0(n1794), .Y(n2511) );
  MXI2X1 U3045 ( .A(n2499), .B(n2495), .S0(n1788), .Y(n2496) );
  INVX1 U3046 ( .A(n2497), .Y(n2494) );
  INVX1 U3047 ( .A(n2506), .Y(n2491) );
  INVX1 U3048 ( .A(n2505), .Y(n2492) );
  NOR2X1 U3049 ( .A(n2519), .B(n2504), .Y(n2505) );
  MXI2X1 U3050 ( .A(n2501), .B(n2500), .S0(n1788), .Y(n2512) );
  INVX1 U3051 ( .A(n2499), .Y(n2500) );
  AND3X1 U3052 ( .A(n2529), .B(n2528), .C(n2701), .Y(n2497) );
  INVX1 U3053 ( .A(n2504), .Y(n2701) );
  MXI2X2 U3054 ( .A(n2560), .B(n2559), .S0(n995), .Y(n2721) );
  INVX1 U3055 ( .A(n2558), .Y(n2559) );
  MXI2X1 U3056 ( .A(n2646), .B(n2645), .S0(n1794), .Y(n2551) );
  AOI2BB2X1 U3057 ( .B0(n2550), .B1(n2694), .A0N(n1265), .A1N(n2549), .Y(n2647) );
  INVX1 U3058 ( .A(n2667), .Y(n2549) );
  INVX1 U3059 ( .A(n2557), .Y(n2560) );
  MXI2X1 U3060 ( .A(n2645), .B(n2646), .S0(n1794), .Y(n2552) );
  MXI2X1 U3061 ( .A(n2541), .B(n2540), .S0(n1788), .Y(n2646) );
  MXI2X1 U3062 ( .A(n2547), .B(n2548), .S0(n1008), .Y(n2645) );
  INVX1 U3063 ( .A(n2546), .Y(n2527) );
  MXI2X1 U3064 ( .A(n2543), .B(n2542), .S0(n1788), .Y(n2553) );
  INVX1 U3065 ( .A(n2541), .Y(n2542) );
  INVX1 U3066 ( .A(n2540), .Y(n2543) );
  INVX1 U3067 ( .A(n2529), .Y(n2530) );
  INVX1 U3068 ( .A(n2528), .Y(n2531) );
  INVX1 U3069 ( .A(n2532), .Y(n2533) );
  MXI2X2 U3070 ( .A(n2556), .B(n2555), .S0(n995), .Y(n2720) );
  INVX1 U3071 ( .A(n2571), .Y(n2555) );
  INVX1 U3072 ( .A(n2570), .Y(n2556) );
  INVX1 U3073 ( .A(n2737), .Y(n2671) );
  MXI2X1 U3074 ( .A(n2572), .B(n1120), .S0(n998), .Y(n2737) );
  INVX1 U3075 ( .A(n2525), .Y(n2516) );
  INVX1 U3076 ( .A(n2524), .Y(n2517) );
  MXI2X1 U3077 ( .A(n2525), .B(n2524), .S0(n1796), .Y(n2570) );
  MXI2X1 U3078 ( .A(n2522), .B(n2523), .S0(n1794), .Y(n2524) );
  NOR2X1 U3079 ( .A(n1788), .B(n2515), .Y(n2525) );
  INVX1 U3080 ( .A(n2514), .Y(n2515) );
  MXI2X1 U3081 ( .A(n2566), .B(n2565), .S0(n1780), .Y(n2571) );
  MXI2X1 U3082 ( .A(n2523), .B(n2522), .S0(n1794), .Y(n2565) );
  NAND2X1 U3083 ( .A(n1788), .B(n2514), .Y(n2523) );
  AOI2BB2X1 U3084 ( .B0(n2550), .B1(n2698), .A0N(n1265), .A1N(n2575), .Y(n2566) );
  INVX1 U3085 ( .A(n2519), .Y(n2520) );
  INVX1 U3086 ( .A(n2518), .Y(n2521) );
  INVX1 U3087 ( .A(n1058), .Y(n2698) );
  NOR2X1 U3088 ( .A(n1798), .B(n2860), .Y(n2550) );
  NAND2X1 U3089 ( .A(n1815), .B(n2926), .Y(n821) );
  NAND2BX1 U3090 ( .AN(n3054), .B(n2932), .Y(n733) );
  NAND2BX1 U3091 ( .AN(n3051), .B(n2932), .Y(n738) );
  NAND2X1 U3092 ( .A(n1727), .B(n2932), .Y(n783) );
  NAND2X1 U3093 ( .A(n1721), .B(n2932), .Y(n723) );
  NAND2X1 U3094 ( .A(n2938), .B(n1713), .Y(n772) );
  NAND2X1 U3095 ( .A(n2938), .B(n1731), .Y(n771) );
  NAND2X1 U3096 ( .A(n2938), .B(n3068), .Y(n2641) );
  AOI2BB2X1 U3097 ( .B0(tree_mem[1]), .B1(n2924), .A0N(tree_mem[1]), .A1N(
        n2924), .Y(n823) );
  NOR2X1 U3098 ( .A(n1715), .B(n2921), .Y(n2924) );
  NAND2X1 U3099 ( .A(n2925), .B(n1702), .Y(n2921) );
  NAND2X1 U3100 ( .A(n2938), .B(n2931), .Y(n784) );
  NAND2X1 U3101 ( .A(n2934), .B(n1716), .Y(n780) );
  NAND2X1 U3102 ( .A(n1722), .B(n2934), .Y(n779) );
  NAND2X1 U3103 ( .A(n1730), .B(n2934), .Y(n778) );
  NAND2BX1 U3104 ( .AN(out_en), .B(n2930), .Y(n762) );
  NAND2BX1 U3105 ( .AN(n2920), .B(n1732), .Y(n825) );
  NAND2X1 U3106 ( .A(n1701), .B(n2930), .Y(n756) );
  NAND2X1 U3107 ( .A(n1693), .B(n2930), .Y(n763) );
  NAND2BX1 U3108 ( .AN(n2927), .B(n2912), .Y(n2926) );
  AOI2BB2X1 U3109 ( .B0(n2934), .B1(n3065), .A0N(n2642), .A1N(n1733), .Y(n2643) );
  OAI2BB1X1 U3110 ( .A0N(n810), .A1N(n2582), .B0(n2913), .Y(n2642) );
  NAND2X1 U3111 ( .A(n2929), .B(n2930), .Y(n2928) );
  OAI2BB1X1 U3112 ( .A0N(n3070), .A1N(n2910), .B0(n2941), .Y(n768) );
  OAI2BB1X1 U3113 ( .A0N(n3071), .A1N(n2910), .B0(n2941), .Y(n707) );
  OAI2BB1X1 U3114 ( .A0N(n3067), .A1N(n2910), .B0(n2940), .Y(n769) );
  OAI2BB1X1 U3115 ( .A0N(n3066), .A1N(n2910), .B0(n2940), .Y(n708) );
  INVX1 U3116 ( .A(n2936), .Y(n2583) );
  NAND2X1 U3117 ( .A(n1741), .B(n2939), .Y(n2950) );
  AOI2BB2X1 U3118 ( .B0(n1814), .B1(n529), .A0N(n1814), .A1N(n3100), .Y(n729)
         );
  AOI2BB2X1 U3119 ( .B0(n1814), .B1(n553), .A0N(n1814), .A1N(n3078), .Y(n742)
         );
  AOI2BB2X1 U3120 ( .B0(n1814), .B1(n475), .A0N(n1814), .A1N(n3107), .Y(n699)
         );
  NAND2X1 U3121 ( .A(n474), .B(n1814), .Y(n698) );
  AOI2BB2X1 U3122 ( .B0(n1814), .B1(n507), .A0N(n1814), .A1N(n3090), .Y(n717)
         );
  AOI2BB2X1 U3123 ( .B0(n1814), .B1(n493), .A0N(n1814), .A1N(n3105), .Y(n710)
         );
  AOI2BB2X1 U3124 ( .B0(n1814), .B1(n497), .A0N(n1814), .A1N(n3103), .Y(n712)
         );
  AOI2BB2X1 U3125 ( .B0(n1814), .B1(n505), .A0N(n1814), .A1N(n3091), .Y(n716)
         );
  AOI2BB2X1 U3126 ( .B0(n1814), .B1(n509), .A0N(n1814), .A1N(n3089), .Y(n718)
         );
  AOI2BB2X1 U3127 ( .B0(n1814), .B1(n524), .A0N(n1814), .A1N(n3086), .Y(n726)
         );
  AOI2BB2X1 U3128 ( .B0(n1814), .B1(n522), .A0N(n1814), .A1N(n3096), .Y(n725)
         );
  AOI2BB2X1 U3129 ( .B0(n1814), .B1(n511), .A0N(n1814), .A1N(n3088), .Y(n719)
         );
  AOI2BB2X1 U3130 ( .B0(n1814), .B1(n520), .A0N(n1814), .A1N(n3101), .Y(n724)
         );
  AOI2BB2X1 U3131 ( .B0(n1814), .B1(n491), .A0N(n1814), .A1N(n3106), .Y(n709)
         );
  AOI2BB2X1 U3132 ( .B0(n1814), .B1(n485), .A0N(n1814), .A1N(n3082), .Y(n704)
         );
  AOI2BB2X1 U3133 ( .B0(n1814), .B1(n483), .A0N(n1814), .A1N(n3087), .Y(n703)
         );
  AOI2BB2X1 U3134 ( .B0(n1814), .B1(n477), .A0N(n1814), .A1N(n3102), .Y(n700)
         );
  AOI2BB2X1 U3135 ( .B0(n1814), .B1(n551), .A0N(n1814), .A1N(n3083), .Y(n741)
         );
  AOI2BB2X1 U3136 ( .B0(n1814), .B1(n526), .A0N(n1814), .A1N(n3081), .Y(n727)
         );
  AOI2BB2X1 U3137 ( .B0(n1814), .B1(n544), .A0N(n1814), .A1N(n3079), .Y(n737)
         );
  AOI2BB2X1 U3138 ( .B0(n1814), .B1(n495), .A0N(n1814), .A1N(n3104), .Y(n711)
         );
  AOI2BB2X1 U3139 ( .B0(n1814), .B1(n549), .A0N(n1814), .A1N(n3093), .Y(n740)
         );
  AOI2BB2X1 U3140 ( .B0(n1814), .B1(n479), .A0N(n1814), .A1N(n3097), .Y(n701)
         );
  AOI2BB2X1 U3141 ( .B0(n1814), .B1(n481), .A0N(n1814), .A1N(n3092), .Y(n702)
         );
  AOI2BB2X1 U3142 ( .B0(n1814), .B1(n547), .A0N(n1814), .A1N(n3098), .Y(n739)
         );
  AOI2BB2X1 U3143 ( .B0(n1814), .B1(n542), .A0N(n1814), .A1N(n3084), .Y(n736)
         );
  OR4X1 U3144 ( .A(gray_valid), .B(n1712), .C(state[1]), .D(state[2]), .Y(
        n2944) );
  NAND2X1 U3145 ( .A(n1783), .B(N774), .Y(n1843) );
  NAND2X1 U3146 ( .A(n1783), .B(N781), .Y(n1844) );
  NAND2X1 U3147 ( .A(n1875), .B(N810), .Y(n1869) );
  NAND2X1 U3148 ( .A(n1875), .B(N809), .Y(n1870) );
  NAND2X1 U3149 ( .A(n1875), .B(N812), .Y(n1867) );
  NAND2X1 U3150 ( .A(n1875), .B(N806), .Y(n1873) );
  NAND2X1 U3151 ( .A(n1875), .B(N807), .Y(n1872) );
  NAND2X1 U3152 ( .A(n1875), .B(N813), .Y(n1874) );
  NAND2X1 U3153 ( .A(n1875), .B(N808), .Y(n1871) );
  NAND2X1 U3154 ( .A(n1875), .B(N811), .Y(n1868) );
  NAND2X1 U3155 ( .A(n1783), .B(N778), .Y(n1839) );
  NAND2X1 U3156 ( .A(n1783), .B(N777), .Y(n1840) );
  NAND2X1 U3157 ( .A(n1783), .B(N775), .Y(n1842) );
  NAND2X1 U3158 ( .A(n1783), .B(N779), .Y(n1838) );
  NAND2X1 U3159 ( .A(n1783), .B(N780), .Y(n1837) );
  NAND2X1 U3160 ( .A(n1783), .B(N776), .Y(n1841) );
  NAND2X1 U3161 ( .A(n1782), .B(N790), .Y(n1825) );
  NAND2X1 U3162 ( .A(n1782), .B(N797), .Y(n1826) );
  NAND2X1 U3163 ( .A(n1782), .B(N792), .Y(n1823) );
  NAND2X1 U3164 ( .A(n1782), .B(N796), .Y(n1819) );
  NAND2X1 U3165 ( .A(n1782), .B(N794), .Y(n1821) );
  NAND2X1 U3166 ( .A(n1782), .B(N795), .Y(n1820) );
  NAND2X1 U3167 ( .A(n1782), .B(N793), .Y(n1822) );
  NAND2X1 U3168 ( .A(n1782), .B(N791), .Y(n1824) );
  NAND2X1 U3169 ( .A(n1836), .B(N770), .Y(n1830) );
  NAND2X1 U3170 ( .A(n1836), .B(N768), .Y(n1832) );
  NAND2X1 U3171 ( .A(n1855), .B(N782), .Y(n1853) );
  NAND2X1 U3172 ( .A(n1836), .B(N767), .Y(n1833) );
  NAND2X1 U3173 ( .A(n1836), .B(N769), .Y(n1831) );
  NAND2X1 U3174 ( .A(n1836), .B(N766), .Y(n1834) );
  NAND2X1 U3175 ( .A(n1855), .B(N786), .Y(n1849) );
  NAND2X1 U3176 ( .A(n1855), .B(N788), .Y(n1847) );
  NAND2X1 U3177 ( .A(n1855), .B(N785), .Y(n1850) );
  NAND2X1 U3178 ( .A(n1836), .B(N771), .Y(n1829) );
  NAND2X1 U3179 ( .A(n1855), .B(N789), .Y(n1854) );
  NAND2X1 U3180 ( .A(n1836), .B(N773), .Y(n1835) );
  NAND2X1 U3181 ( .A(n1836), .B(N772), .Y(n1828) );
  NAND2X1 U3182 ( .A(n1855), .B(N784), .Y(n1851) );
  NAND2X1 U3183 ( .A(n1855), .B(N787), .Y(n1848) );
  NAND2X1 U3184 ( .A(n1855), .B(N783), .Y(n1852) );
  NAND2X1 U3185 ( .A(n1864), .B(N801), .Y(n1859) );
  NAND2X1 U3186 ( .A(n1864), .B(N802), .Y(n1858) );
  NAND2X1 U3187 ( .A(n1864), .B(N803), .Y(n1857) );
  NAND2X1 U3188 ( .A(n1864), .B(N799), .Y(n1861) );
  NAND2X1 U3189 ( .A(n1864), .B(N805), .Y(n1863) );
  NAND2X1 U3190 ( .A(n1864), .B(N800), .Y(n1860) );
  NAND2X1 U3191 ( .A(n1864), .B(N804), .Y(n1856) );
  NAND2X1 U3192 ( .A(n1864), .B(N798), .Y(n1862) );
  NAND3X1 U3193 ( .A(gray_data[1]), .B(gray_data[0]), .C(gray_data[2]), .Y(
        n2919) );
  NOR4X1 U3194 ( .A(gray_data[7]), .B(gray_data[6]), .C(gray_data[5]), .D(
        gray_data[4]), .Y(n2918) );
  NAND2BX1 U3195 ( .AN(n629), .B(n2282), .Y(n2278) );
  NAND2BX1 U3196 ( .AN(n630), .B(n2282), .Y(n2277) );
  NAND2BX1 U3197 ( .AN(n631), .B(n2282), .Y(n2276) );
  NAND2BX1 U3198 ( .AN(n632), .B(n2282), .Y(n2281) );
  NAND2BX1 U3199 ( .AN(n633), .B(n2282), .Y(n2280) );
  NAND2BX1 U3200 ( .AN(n634), .B(n2282), .Y(n2274) );
  NAND2BX1 U3201 ( .AN(n635), .B(n2282), .Y(n2272) );
  NAND2BX1 U3202 ( .AN(n636), .B(n2282), .Y(n2283) );
  NOR2X1 U3203 ( .A(n2332), .B(n2438), .Y(n2323) );
  OAI21X1 U3204 ( .A0(n2772), .A1(n2910), .B0(n2771), .Y(n706) );
  NAND2X1 U3205 ( .A(n2910), .B(n3076), .Y(n2771) );
  AOI211X1 U3206 ( .A0(n2763), .A1(\com[0][4] ), .B0(n2762), .C0(n2761), .Y(
        n2764) );
  INVX1 U3207 ( .A(\com[1][2] ), .Y(n2756) );
  INVX1 U3208 ( .A(\com[0][0] ), .Y(n2751) );
  INVX1 U3209 ( .A(\com[0][1] ), .Y(n2752) );
  INVX1 U3210 ( .A(\com[1][4] ), .Y(n2763) );
  INVX1 U3211 ( .A(n2761), .Y(n2766) );
  INVX1 U3212 ( .A(\com[0][5] ), .Y(n2750) );
  INVX1 U3213 ( .A(\com[0][6] ), .Y(n2768) );
  NAND2BX1 U3214 ( .AN(n613), .B(n2448), .Y(n2439) );
  NAND2X1 U3215 ( .A(\com[3][5] ), .B(n623), .Y(n2376) );
  OAI211X1 U3216 ( .A0(n2485), .A1(n818), .B0(n2484), .C0(n2483), .Y(n2486) );
  INVX1 U3217 ( .A(n2935), .Y(n2483) );
  NAND2X1 U3218 ( .A(n2936), .B(tree_mem_back[0]), .Y(n2935) );
  OAI2BB1X1 U3219 ( .A0N(n2482), .A1N(n2481), .B0(n2480), .Y(n2488) );
  INVX1 U3220 ( .A(n2937), .Y(n2474) );
  NAND2X1 U3221 ( .A(n2936), .B(n1734), .Y(n2937) );
  NOR2X1 U3222 ( .A(n2345), .B(n622), .Y(n2346) );
  AOI21X1 U3223 ( .A0(n2345), .A1(n622), .B0(com_after_1[6]), .Y(n2347) );
  AOI21X1 U3224 ( .A0(n2342), .A1(n2341), .B0(n2340), .Y(n2344) );
  NOR2X1 U3226 ( .A(n2337), .B(n2336), .Y(n2339) );
  NOR2X1 U3227 ( .A(n629), .B(n809), .Y(n2337) );
  INVX1 U3228 ( .A(n2932), .Y(n2350) );
  INVX1 U3229 ( .A(n2629), .Y(n2625) );
  INVX1 U3230 ( .A(n2633), .Y(n2621) );
  NAND2X1 U3231 ( .A(n2948), .B(n605), .Y(n2629) );
  NOR2X1 U3232 ( .A(n2929), .B(n1729), .Y(n2948) );
  INVX1 U3233 ( .A(n2938), .Y(n2454) );
  NAND2BX1 U3234 ( .AN(n608), .B(n2592), .Y(n2591) );
  INVX1 U3235 ( .A(n1953), .Y(n1966) );
  MXI2X1 U3236 ( .A(n1214), .B(n1203), .S0(n1325), .Y(n1953) );
  AND2X1 U3237 ( .A(n2987), .B(n2690), .Y(n1754) );
  AO22X1 U3238 ( .A0(n2957), .A1(n2958), .B0(n2906), .B1(n2959), .Y(n2956) );
  OA22X1 U3239 ( .A0(n2849), .A1(n1708), .B0(n2850), .B1(n1697), .Y(n1751) );
  OA22X1 U3240 ( .A0(n2849), .A1(n1709), .B0(n2850), .B1(n1698), .Y(n1752) );
  OA22X1 U3241 ( .A0(n2853), .A1(n1708), .B0(n2854), .B1(n1697), .Y(n1748) );
  OA22X1 U3242 ( .A0(n2853), .A1(n1709), .B0(n2854), .B1(n1698), .Y(n1749) );
  OA22X1 U3243 ( .A0(n2853), .A1(n1705), .B0(n2854), .B1(n1118), .Y(n1744) );
  OA22X1 U3244 ( .A0(n2853), .A1(n1706), .B0(n2854), .B1(n1696), .Y(n1745) );
  OA22X1 U3245 ( .A0(n2853), .A1(n1699), .B0(n2854), .B1(n1707), .Y(n1750) );
  OA22X1 U3246 ( .A0(n2849), .A1(n1706), .B0(n2850), .B1(n1696), .Y(n1747) );
  OA22X1 U3247 ( .A0(n2849), .A1(n1699), .B0(n2850), .B1(n1707), .Y(n1753) );
  AND4X1 U3248 ( .A(n2739), .B(n2738), .C(n2788), .D(n2737), .Y(n2777) );
  OAI21XL U3249 ( .A0(n1734), .A1(n2929), .B0(tree_mem_back[1]), .Y(n2931) );
  NOR2BX1 U3257 ( .AN(n2916), .B(gray_data[0]), .Y(n1827) );
  OAI21XL U3258 ( .A0(n2692), .A1(n2745), .B0(n2957), .Y(n3000) );
  OAI31XL U3259 ( .A0(n2777), .A1(n2806), .A2(n2748), .B0(n2747), .Y(n2749) );
  OAI31XL U3260 ( .A0(n2802), .A1(n2736), .A2(n2801), .B0(n2554), .Y(n2955) );
  OAI22XL U3261 ( .A0(n1701), .A1(n2852), .B0(n2828), .B1(n1721), .Y(n3011) );
  OAI22XL U3262 ( .A0(n2859), .A1(n1705), .B0(n2860), .B1(n1118), .Y(n2836) );
  OA21XL U3263 ( .A0(n1731), .A1(n2824), .B0(n2658), .Y(n2953) );
  OAI22XL U3264 ( .A0(n1693), .A1(n2859), .B0(n2860), .B1(n1701), .Y(n2656) );
  OA21XL U3265 ( .A0(n1721), .A1(n2827), .B0(n2726), .Y(n3026) );
  OAI22XL U3266 ( .A0(n1701), .A1(n2856), .B0(n1693), .B1(n2855), .Y(n2970) );
  OAI22XL U3267 ( .A0(n1693), .A1(n2853), .B0(n1701), .B1(n2854), .Y(n2993) );
  OAI22XL U3268 ( .A0(n2854), .A1(n1695), .B0(n1704), .B1(n2853), .Y(n2812) );
  OR2X1 U3269 ( .A(n2908), .B(n2680), .Y(n2682) );
  OAI22XL U3270 ( .A0(n2859), .A1(n1706), .B0(n2860), .B1(n1696), .Y(n2833) );
  OAI22XL U3271 ( .A0(n1704), .A1(n2855), .B0(n1695), .B1(n2856), .Y(n2817) );
  OAI21XL U3272 ( .A0(n2736), .A1(n2801), .B0(n2986), .Y(n2984) );
  OAI22XL U3273 ( .A0(n2850), .A1(n1695), .B0(n1704), .B1(n2849), .Y(n2790) );
  OA21XL U3274 ( .A0(n2801), .A1(n2959), .B0(n2906), .Y(n2789) );
  OAI22XL U3275 ( .A0(n2852), .A1(n1695), .B0(n2851), .B1(n1704), .Y(n2807) );
  OAI21XL U3276 ( .A0(n2736), .A1(n2906), .B0(n2959), .Y(n2738) );
  OAI22XL U3277 ( .A0(n2848), .A1(n1704), .B0(n2847), .B1(n1695), .Y(n2773) );
  OA21XL U3278 ( .A0(n2733), .A1(n2981), .B0(n2747), .Y(n2776) );
  OAI222XL U3279 ( .A0(n1097), .A1(n2847), .B0(n1694), .B1(n3040), .C0(n2848), 
        .C1(n1114), .Y(N648) );
  OAI22XL U3280 ( .A0(n2901), .A1(n2716), .B0(n2712), .B1(n2711), .Y(n2717) );
  OR2X1 U3281 ( .A(n1058), .B(n2701), .Y(n2702) );
  OAI22XL U3282 ( .A0(n2860), .A1(n1695), .B0(n2859), .B1(n1704), .Y(n2822) );
  OR2X1 U3283 ( .A(n2683), .B(n2654), .Y(n2655) );
  OAI21XL U3284 ( .A0(n2674), .A1(n2649), .B0(n2652), .Y(n2654) );
  AND2X1 U3285 ( .A(n3045), .B(n3020), .Y(n1743) );
  OAI21XL U3286 ( .A0(n2529), .A1(n2493), .B0(n2528), .Y(n2499) );
  NAND2XL U3287 ( .A(tree_mem_back[1]), .B(n775), .Y(n2473) );
  AOI211XL U3288 ( .A0(state[1]), .A1(n2945), .B0(n2946), .C0(state[2]), .Y(
        n2943) );
  NAND3XL U3289 ( .A(n3108), .B(n2912), .C(n1712), .Y(n2945) );
  OAI22XL U3290 ( .A0(n2753), .A1(\com[1][2] ), .B0(\com[1][1] ), .B1(n2752), 
        .Y(n2754) );
  OAI22XL U3291 ( .A0(com_after_1[5]), .A1(n623), .B0(n624), .B1(
        com_after_1[4]), .Y(n2343) );
  OAI22XL U3292 ( .A0(n806), .A1(n632), .B0(n633), .B1(n805), .Y(n2340) );
  OAI22XL U3293 ( .A0(n2339), .A1(n2338), .B0(n807), .B1(n631), .Y(n2342) );
  OAI22XL U3294 ( .A0(com_after_1[2]), .A1(n626), .B0(n627), .B1(
        com_after_1[1]), .Y(n2338) );
  OR2X1 U3295 ( .A(n2948), .B(n2865), .Y(n2633) );
  OAI21XL U3296 ( .A0(n2600), .A1(n792), .B0(n2599), .Y(n2606) );
  OR2X1 U3297 ( .A(n2938), .B(n613), .Y(n1700) );
  OR2X1 U3298 ( .A(tree_mem_back[1]), .B(tree_mem_back[0]), .Y(n1729) );
  AO21X1 U3299 ( .A0(tree_mem[0]), .A1(n2921), .B0(n2922), .Y(n824) );
  OAI31XL U3300 ( .A0(n1736), .A1(n2923), .A2(n1715), .B0(n1702), .Y(n822) );
  OAI31XL U3301 ( .A0(n1720), .A1(n2927), .A2(n1738), .B0(n1740), .Y(n819) );
  OAI21XL U3302 ( .A0(n2913), .A1(n1718), .B0(n2933), .Y(n781) );
  OAI21XL U3303 ( .A0(n2911), .A1(n1703), .B0(n2942), .Y(n767) );
  OR2X1 U3304 ( .A(n3053), .B(n2911), .Y(n766) );
  OR2X1 U3305 ( .A(n3056), .B(n2911), .Y(n765) );
  OR2X1 U3306 ( .A(n3059), .B(n2911), .Y(n764) );
  OAI22XL U3307 ( .A0(n2920), .A1(n1737), .B0(n1740), .B1(n2926), .Y(n761) );
  OAI21XL U3308 ( .A0(n2911), .A1(n1115), .B0(n2942), .Y(n760) );
  OR2X1 U3309 ( .A(n3052), .B(n2911), .Y(n759) );
  OR2X1 U3310 ( .A(n3055), .B(n2911), .Y(n758) );
  OR2X1 U3311 ( .A(n3060), .B(n2911), .Y(n757) );
  OR2X1 U3312 ( .A(n2948), .B(n3061), .Y(n705) );
  OAI21XL U3313 ( .A0(n1114), .A1(n2939), .B0(n2949), .Y(n695) );
  OAI21XL U3314 ( .A0(n1097), .A1(n2939), .B0(n2949), .Y(n694) );
  OAI221XL U3315 ( .A0(tree_mem_back[1]), .A1(n3064), .B0(n1741), .B1(n3068), 
        .C0(n2939), .Y(n2949) );
  OAI222XL U3316 ( .A0(n1694), .A1(n2936), .B0(n2937), .B1(n1733), .C0(n1717), 
        .C1(n2935), .Y(n692) );
  OAI22XL U3317 ( .A0(n1694), .A1(n2950), .B0(n2939), .B1(n1113), .Y(n691) );
  OAI22XL U3318 ( .A0(n1694), .A1(n2950), .B0(n2939), .B1(n1096), .Y(n690) );
  OAI21XL U3319 ( .A0(n2966), .A1(n1731), .B0(n2969), .Y(N706) );
  OAI22XL U3320 ( .A0(n2961), .A1(n1730), .B0(n1723), .B1(n2972), .Y(n2971) );
  OAI21XL U3321 ( .A0(n2904), .A1(n2981), .B0(n2982), .Y(n2980) );
  OAI21XL U3322 ( .A0(n1730), .A1(n2987), .B0(n2992), .Y(N692) );
  OAI22XL U3323 ( .A0(n1731), .A1(n2991), .B0(n1723), .B1(n2995), .Y(n2994) );
  OAI21XL U3324 ( .A0(n1730), .A1(n3002), .B0(n3010), .Y(N678) );
  OAI22XL U3325 ( .A0(n1731), .A1(n3009), .B0(n1723), .B1(n3013), .Y(n3012) );
  OAI21XL U3326 ( .A0(n1730), .A1(n3021), .B0(n3026), .Y(N664) );
  OAI22XL U3327 ( .A0(n1731), .A1(n3025), .B0(n1723), .B1(n3028), .Y(n3027) );
  OAI21XL U3328 ( .A0(n3031), .A1(n1730), .B0(n3039), .Y(N650) );
  OAI21XL U3329 ( .A0(n1732), .A1(n2923), .B0(n2951), .Y(N205) );
  OAI221XL U3330 ( .A0(state[2]), .A1(gray_valid), .B0(n1711), .B1(out_en), 
        .C0(n1725), .Y(n3048) );
  OAI221XL U3331 ( .A0(state[0]), .A1(n3077), .B0(n1712), .B1(n1732), .C0(
        state[1]), .Y(n3047) );
  huffman_DW01_inc_0 add_227 ( .A(CNT6), .SUM({N813, N812, N811, N810, N809, 
        N808, N807, N806}) );
  huffman_DW01_inc_1 add_224 ( .A(CNT5), .SUM({N805, N804, N803, N802, N801, 
        N800, N799, N798}) );
  huffman_DW01_inc_2 add_221 ( .A(CNT4), .SUM({N797, N796, N795, N794, N793, 
        N792, N791, N790}) );
  huffman_DW01_inc_3 add_218 ( .A(CNT3), .SUM({N789, N788, N787, N786, N785, 
        N784, N783, N782}) );
  huffman_DW01_inc_4 add_215 ( .A({n1196, CNT2[6:0]}), .SUM({N781, N780, N779, 
        N778, N777, N776, N775, N774}) );
  huffman_DW01_inc_5 add_212 ( .A({CNT1[7:5], n1204, CNT1[3:0]}), .SUM({N773, 
        N772, N771, N770, N769, N768, N767, N766}) );
  huffman_DW01_add_2 add_323 ( .A({n794, n795, n796, n797, n798, n799, n800, 
        n801}), .B({1'b0, \com[4][6] , \com[4][5] , \com[4][4] , \com[4][3] , 
        \com[4][2] , \com[4][1] , \com[4][0] }), .CI(1'b0), .SUM({N1222, N1221, 
        N1220, N1219, N1218, N1217, N1216, N1215}), .IN0(clk), .IN1(n1813), 
        .IN2(n1809), .IN3(n1808), .IN4(n3123) );
  huffman_add_314_DP_OP_292_9816_0 add_314_DP_OP_292_9816_3 ( .I1({n818, 
        com_after_1[6:0]}), .I2({n802, n803, n804, n805, n806, n807, n808, 
        n809}), .O2({n2897, n2896, n2895, n2894, n2893, n2892, n2891, n2890})
         );
  huffman_add_318_DP_OP_291_9816_1 add_318_DP_OP_291_9816_4 ( .I1({n802, n803, 
        n804, n805, n806, n807, n808, n809}), .I2({\com[3][7] , \com[3][6] , 
        \com[3][5] , \com[3][4] , \com[3][3] , n1100, \com[3][1] , \com[3][0] }), .O1({n2889, n2888, n2887, n2886, n2885, n2884, n2883, n2882}), .IN0(clk), 
        .IN1(n1813), .IN2(n1808) );
  huffman_add_303_DP_OP_294_9816_1 add_303_DP_OP_294_9816_5 ( .I1({\com[3][7] , 
        \com[3][6] , \com[3][5] , \com[3][4] , \com[3][3] , n1100, \com[3][1] , 
        \com[3][0] }), .I2({\com[2][7] , \com[2][6] , \com[2][5] , \com[2][4] , 
        \com[2][3] , \com[2][2] , \com[2][1] , \com[2][0] }), .O2({n2881, 
        n2880, n2879, n2878, n2877, n2876, n2875, n2874}), .IN0(clk), .IN1(
        n1813), .IN2(n1808), .IN3(n1809) );
  huffman_add_307_DP_OP_293_9816_1 add_307_DP_OP_293_9816_6 ( .I1({n818, 
        com_after_1[6:0]}), .I2({\com[2][7] , \com[2][6] , \com[2][5] , 
        \com[2][4] , \com[2][3] , \com[2][2] , \com[2][1] , \com[2][0] }), 
        .O1({n2873, n2872, n2871, n2870, n2869, n2868, n2867, n2866}) );
  huffman_DW01_add_13 add_297 ( .A({\com[0][7] , \com[0][6] , \com[0][5] , 
        \com[0][4] , \com[0][3] , \com[0][2] , \com[0][1] , \com[0][0] }), .B(
        {\com[1][7] , \com[1][6] , n1191, \com[1][4] , \com[1][3] , 
        \com[1][2] , \com[1][1] , \com[1][0] }), .CI(1'b0), .SUM({N1147, N1146, 
        N1145, N1144, N1143, N1142, N1141, N1140}) );
  DFFSX1 R_2 ( .D(n2590), .CK(clk), .SN(n1813), .Q(n3254) );
  DFFSX1 R_5 ( .D(n2593), .CK(clk), .SN(n1809), .Q(n3253) );
  DFFSXL R_8 ( .D(n2589), .CK(clk), .SN(n1808), .Q(n3252) );
  DFFSXL R_9 ( .D(n2592), .CK(clk), .SN(n1813), .Q(n3251) );
  DFFSX1 R_17 ( .D(n2591), .CK(clk), .SN(n1813), .Q(n3250) );
  MXI2X4 U1779 ( .A(n2326), .B(n3249), .S0(n3127), .Y(n805) );
  DFFSX1 R_26 ( .D(n624), .CK(clk), .SN(n1809), .Q(n3249) );
  DFFSX1 R_35 ( .D(n610), .CK(clk), .SN(n1813), .Q(n3248) );
  DFFSX1 R_38 ( .D(n623), .CK(clk), .SN(n1813), .Q(n3247) );
  DFFSXL R_43 ( .D(n627), .CK(clk), .SN(n1808), .Q(n3246) );
  DFFSX1 R_46 ( .D(n626), .CK(clk), .SN(n1810), .Q(n3245) );
  DFFSX1 R_52 ( .D(n628), .CK(clk), .SN(n1808), .Q(n3243) );
  NAND2X1 U2583 ( .A(n3170), .B(n3122), .Y(n2458) );
  DFFSXL R_57 ( .D(n617), .CK(clk), .SN(n1813), .Q(n3242) );
  DFFSXL R_60 ( .D(n614), .CK(clk), .SN(n1813), .Q(n3241) );
  DFFSXL R_63 ( .D(n619), .CK(clk), .SN(n1813), .Q(n3240) );
  DFFRX1 R_75 ( .D(n1095), .CK(clk), .RN(n1813), .Q(n3239) );
  DFFSX1 R_76 ( .D(n2913), .CK(clk), .SN(n1813), .Q(n3238) );
  DFFSX1 R_77 ( .D(n1116), .CK(clk), .SN(n1813), .Q(n3237) );
  DFFSX1 R_79 ( .D(n620), .CK(clk), .SN(n1813), .Q(n3236) );
  DFFSX1 R_86 ( .D(n2439), .CK(clk), .SN(n1813), .Q(n3235) );
  DFFSX1 R_90 ( .D(n2936), .CK(clk), .SN(n1813), .Q(n3234) );
  DFFSX1 R_91 ( .D(n1735), .CK(clk), .SN(n1813), .Q(n3233) );
  DFFSX1 R_93 ( .D(n2489), .CK(clk), .SN(n1813), .Q(n3232) );
  OAI22X1 U2439 ( .A0(n2367), .A1(n807), .B0(n2371), .B1(n806), .Y(n2368) );
  DFFSX1 R_98 ( .D(n1135), .CK(clk), .SN(n1809), .Q(n3230) );
  DFFSX1 R_100 ( .D(n1056), .CK(clk), .SN(n1813), .Q(n3229) );
  DFFSX1 R_104 ( .D(n2582), .CK(clk), .SN(n1813), .Q(n3228) );
  DFFSX1 R_105 ( .D(n1692), .CK(clk), .SN(n1813), .Q(n3227) );
  DFFSX1 R_111 ( .D(n2625), .CK(clk), .SN(n1812), .Q(n3226) );
  DFFSX1 R_127 ( .D(n616), .CK(clk), .SN(n1813), .Q(n3225) );
  DFFSX1 R_130 ( .D(n612), .CK(clk), .SN(n1813), .Q(n3224) );
  DFFRX1 R_133 ( .D(n2871), .CK(clk), .RN(n1813), .Q(n3223) );
  DFFRX1 R_136 ( .D(n2870), .CK(clk), .RN(n1809), .Q(n3222) );
  DFFRX1 R_146 ( .D(n2474), .CK(clk), .RN(n1813), .Q(n3220) );
  DFFSX1 R_151 ( .D(n2873), .CK(clk), .SN(n1808), .Q(n3218) );
  DFFSX1 R_154 ( .D(n621), .CK(clk), .SN(n1808), .Q(n3217) );
  DFFSX1 R_155 ( .D(n2876), .CK(clk), .SN(n1810), .Q(n3216) );
  DFFRX1 R_156 ( .D(n2868), .CK(clk), .RN(n1810), .Q(n3215) );
  DFFSX1 R_158 ( .D(n1446), .CK(clk), .SN(n1813), .Q(n3214) );
  DFFSX1 R_162 ( .D(n2874), .CK(clk), .SN(n1808), .Q(n3212) );
  DFFRX1 R_163 ( .D(n2866), .CK(clk), .RN(n1808), .Q(n3211) );
  DFFSX1 R_170 ( .D(n2608), .CK(clk), .SN(n1812), .Q(n3210) );
  DFFSX1 R_171 ( .D(n611), .CK(clk), .SN(n1812), .Q(n3209) );
  DFFSX1 R_181 ( .D(n2631), .CK(clk), .SN(n1812), .Q(n3208) );
  DFFSX1 R_183 ( .D(\com[4][2] ), .CK(clk), .SN(n1813), .Q(n3207) );
  DFFSX1 R_192 ( .D(n2872), .CK(clk), .SN(n1813), .Q(n3205) );
  DFFSX1 R_195 ( .D(n622), .CK(clk), .SN(n1813), .Q(n3204) );
  DFFSX1 R_208 ( .D(n2379), .CK(clk), .SN(n1813), .Q(n3201) );
  DFFRX1 R_209 ( .D(\com[3][7] ), .CK(clk), .RN(n1813), .Q(n3200) );
  DFFRX1 R_210 ( .D(n621), .CK(clk), .RN(n1813), .Q(n3199) );
  DFFRX1 R_212 ( .D(n2629), .CK(clk), .RN(n1812), .Q(n3198) );
  DFFSX1 R_223 ( .D(n976), .CK(clk), .SN(n1813), .Q(n3192) );
  DFFSX1 R_230 ( .D(n2438), .CK(clk), .SN(n1813), .Q(n3191) );
  DFFSX1 R_233 ( .D(n613), .CK(clk), .SN(n1813), .Q(n3189) );
  DFFSX1 R_238 ( .D(\com[3][7] ), .CK(clk), .SN(n1813), .Q(n3188) );
  DFFSX1 R_239 ( .D(n2485), .CK(clk), .SN(n1813), .Q(n3187) );
  DFFSX1 R_241 ( .D(n2875), .CK(clk), .SN(n1808), .Q(n3186) );
  DFFRX1 R_242 ( .D(n2867), .CK(clk), .RN(n1808), .Q(n3185) );
  DFFSX1 R_248 ( .D(n2616), .CK(clk), .SN(n1812), .Q(n3184) );
  DFFSX1 R_264 ( .D(n1700), .CK(clk), .SN(n1813), .Q(n3181) );
  DFFSX1 R_265 ( .D(n2454), .CK(clk), .SN(n1813), .Q(n3180) );
  DFFSX1 R_266 ( .D(n1719), .CK(clk), .SN(n1813), .Q(n3179) );
  DFFSX1 R_150_RW ( .D(n1486), .CK(clk), .SN(n1813), .Q(n3219) );
  DFFRX1 R_268 ( .D(\com[4][0] ), .CK(clk), .RN(n1813), .Q(n3178) );
  DFFSX1 R_282 ( .D(n1726), .CK(clk), .SN(n1808), .Q(n3174) );
  DFFSX1 R_283 ( .D(n2323), .CK(clk), .SN(n1808), .Q(n3173) );
  DFFRX1 R_190_RW ( .D(n2438), .CK(clk), .RN(n1808), .Q(n3206) );
  DFFSX1 R_286 ( .D(n1482), .CK(clk), .SN(n1812), .Q(n3172) );
  DFFSX1 R_300 ( .D(n2457), .CK(clk), .SN(n1813), .Q(n3170) );
  DFFSX1 R_303 ( .D(n2452), .CK(clk), .SN(n1813), .Q(n3169) );
  DFFSX1 R_309 ( .D(n2622), .CK(clk), .SN(n1812), .Q(n3167) );
  DFFRX1 R_310 ( .D(n2948), .CK(clk), .RN(n1812), .Q(n3166) );
  DFFRX1 R_311 ( .D(n2621), .CK(clk), .RN(n1812), .Q(n3165) );
  DFFSX1 R_323 ( .D(n2377), .CK(clk), .SN(n1813), .Q(n3164) );
  DFFRX1 R_324 ( .D(n2376), .CK(clk), .RN(n1813), .Q(n3163) );
  DFFSX1 R_325 ( .D(n1449), .CK(clk), .SN(n1813), .Q(n3162) );
  DFFSX1 R_329 ( .D(n1451), .CK(clk), .SN(n1813), .Q(n3160) );
  DFFSX1 R_330 ( .D(n1107), .CK(clk), .SN(n1813), .Q(n3159) );
  DFFRX1 R_331 ( .D(n1448), .CK(clk), .RN(n1813), .Q(n3158) );
  DFFSX1 R_333 ( .D(n2861), .CK(clk), .SN(n1812), .Q(n3157) );
  DFFSX1 R_334 ( .D(n1453), .CK(clk), .SN(n1812), .Q(n3156) );
  DFFRX1 R_335 ( .D(n2607), .CK(clk), .RN(n1812), .Q(n3155) );
  DFFSX1 R_338 ( .D(n1053), .CK(clk), .SN(n1812), .Q(n3154) );
  DFFSX1 R_339 ( .D(n1052), .CK(clk), .SN(n1812), .Q(n3153) );
  DFFRX1 R_343 ( .D(n2625), .CK(clk), .RN(n1812), .Q(n3152) );
  DFFSX1 R_49 ( .D(n615), .CK(clk), .SN(n1813), .Q(n3244) );
  MXI2X2 U2544 ( .A(n2449), .B(n3242), .S0(n3126), .Y(n798) );
  MXI2X4 U1767 ( .A(n3231), .B(n2325), .S0(n3230), .Y(n806) );
  DFFSX1 R_270 ( .D(n801), .CK(clk), .SN(n1813), .Q(n3177) );
  DFFSX1 R_159 ( .D(n800), .CK(clk), .SN(n1813), .Q(n3213) );
  DFFRX1 R_304 ( .D(n795), .CK(clk), .RN(n1813), .Q(n3168) );
  DFFRX1 R_139 ( .D(n797), .CK(clk), .RN(n1813), .Q(n3221) );
  OAI22X1 U2690 ( .A0(n2378), .A1(n802), .B0(n1449), .B1(n803), .Y(n2379) );
  DFFRX1 R_326 ( .D(n803), .CK(clk), .RN(n1813), .Q(n3161) );
  NAND2BX1 U3225 ( .AN(com_after_1[3]), .B(n806), .Y(n2341) );
  AO22X1 U1804 ( .A0(n2372), .A1(n805), .B0(n2371), .B1(n806), .Y(n2373) );
  DFFSX1 R_96 ( .D(n625), .CK(clk), .SN(n1809), .Q(n3231) );
  DFFSX1 R_346 ( .D(n1141), .CK(clk), .SN(n1808), .Q(n3151) );
  DFFRX1 R_201_RW ( .D(n2882), .CK(clk), .RN(n1808), .Q(n3203) );
  DFFSX1 R_202_RW ( .D(n2890), .CK(clk), .SN(n1808), .Q(n3202) );
  DFFRX1 R_213_RW ( .D(n2883), .CK(clk), .RN(n1808), .Q(n3197) );
  DFFSX1 R_214_RW ( .D(n2891), .CK(clk), .SN(n1808), .Q(n3196) );
  DFFRX1 R_216_RW ( .D(n2884), .CK(clk), .RN(n1808), .Q(n3195) );
  DFFSX1 R_217_RW ( .D(n2892), .CK(clk), .SN(n1808), .Q(n3194) );
  DFFRX1 R_219_RW ( .D(n2869), .CK(clk), .RN(n1808), .Q(n3193) );
  DFFSX1 R_231_RW ( .D(n2897), .CK(clk), .SN(n1808), .Q(n3190) );
  DFFSX1 R_254_RW ( .D(n2896), .CK(clk), .SN(n1808), .Q(n3183) );
  DFFSX1 R_257_RW ( .D(n2893), .CK(clk), .SN(n1808), .Q(n3182) );
  DFFSX1 R_275_RW ( .D(n2895), .CK(clk), .SN(n1808), .Q(n3176) );
  DFFSX1 R_279_RW ( .D(n2894), .CK(clk), .SN(n1808), .Q(n3175) );
  CLKINVX1 U2588 ( .A(n2469), .Y(n2455) );
  DFFRX1 R_297 ( .D(n1488), .CK(clk), .RN(n1813), .Q(n3171) );
  DFFRX1 R_380 ( .D(n796), .CK(clk), .RN(n1813), .Q(n3150) );
  DFFSX1 R_383 ( .D(n797), .CK(clk), .SN(n1813), .Q(n3149) );
  DFFSX1 R_385 ( .D(n796), .CK(clk), .SN(n1813), .Q(n3148) );
  DFFSX1 R_391 ( .D(n2596), .CK(clk), .SN(n1812), .Q(n3147) );
  DFFSX1 R_392 ( .D(n2595), .CK(clk), .SN(n1812), .Q(n3146) );
  DFFSX1 R_393 ( .D(n1352), .CK(clk), .SN(n1812), .Q(n3145) );
  DFFSX1 R_397 ( .D(n1466), .CK(clk), .SN(n1812), .Q(n3144) );
  DFFSX1 R_398 ( .D(n606), .CK(clk), .SN(n1812), .Q(n3143) );
  DFFRX2 R_399 ( .D(n2631), .CK(clk), .RN(n1812), .QN(n2618) );
  DFFSX1 R_403 ( .D(n2461), .CK(clk), .SN(n1813), .Q(n3142) );
  DFFSX1 R_404 ( .D(n799), .CK(clk), .SN(n1813), .Q(n3141) );
  DFFSX1 R_409 ( .D(n1460), .CK(clk), .SN(n1812), .Q(n3140) );
  DFFRX1 R_410 ( .D(\com[4][7] ), .CK(clk), .RN(n1813), .Q(n3139) );
  DFFSX1 R_411 ( .D(n1464), .CK(clk), .SN(n1812), .Q(n3138) );
  DFFSX1 R_412 ( .D(n607), .CK(clk), .SN(n1812), .Q(n3137) );
  DFFRX1 R_416 ( .D(n1457), .CK(clk), .RN(n1812), .Q(n3136) );
  DFFRX1 R_417 ( .D(n2863), .CK(clk), .RN(n1812), .Q(n3135) );
  DFFRX1 R_421 ( .D(n2461), .CK(clk), .RN(n1813), .Q(n3134) );
  DFFRX1 R_423 ( .D(n799), .CK(clk), .RN(n1813), .Q(n3133) );
  DFFSX1 R_424 ( .D(n1445), .CK(clk), .SN(n1813), .Q(n3132) );
  DFFRX1 R_425 ( .D(n619), .CK(clk), .RN(n1813), .Q(n3131) );
  DFFSX1 R_430 ( .D(n2284), .CK(clk), .SN(n1810), .Q(n3130) );
  DFFRX1 R_431 ( .D(N1147), .CK(clk), .RN(n1810), .Q(n3129) );
  DFFSX1 R_432 ( .D(n2283), .CK(clk), .SN(n1810), .Q(n3128) );
  DFFSX1 R_440 ( .D(n2594), .CK(clk), .SN(n1813), .Q(n3125) );
  DFFRX1 R_441 ( .D(n2594), .CK(clk), .RN(n1813), .Q(n3124) );
  DFFSX1 R_442 ( .D(\com[4][7] ), .CK(clk), .SN(n1813), .Q(n3123) );
  DFFRX1 R_443 ( .D(n798), .CK(clk), .RN(n1813), .Q(n3122) );
  DFFSX1 R_446 ( .D(n2467), .CK(clk), .SN(n1813), .Q(n3121) );
  DFFSX1 R_447 ( .D(n2468), .CK(clk), .SN(n1813), .Q(n3120) );
  DFFSX1 R_448 ( .D(n2630), .CK(clk), .SN(n1812), .Q(n3119) );
  DFFSX1 R_449 ( .D(n2332), .CK(clk), .SN(n1813), .Q(n3118) );
  DFFSX1 R_450 ( .D(n790), .CK(clk), .SN(n1812), .Q(n3117) );
  DFFRX1 R_451 ( .D(n790), .CK(clk), .RN(n1812), .Q(n3116) );
  DFFSX1 R_452 ( .D(n618), .CK(clk), .SN(n1813), .Q(n3115) );
  DFFSRX2 \hcode3_reg[1]  ( .D(n774), .CK(clk), .SN(1'b1), .RN(n2914), .QN(
        n1714) );
  DFFSRXL \compare_cnt_reg[2]  ( .D(n819), .CK(clk), .SN(1'b1), .RN(n2914), 
        .Q(n3108), .QN(n1740) );
  DFFSX2 R_438 ( .D(n1781), .CK(clk), .SN(n1813), .Q(n3127) );
  DFFSX2 R_439 ( .D(n2448), .CK(clk), .SN(n1813), .Q(n3126) );
  DFFSRX2 \hcode4_reg[2]  ( .D(n773), .CK(clk), .SN(1'b1), .RN(n2914), .Q(
        n3064) );
  INVX3 U1182 ( .A(reset), .Y(n2914) );
  CLKBUFX6 U1185 ( .A(n1810), .Y(n1809) );
  CLKBUFX4 U1186 ( .A(n2914), .Y(n1810) );
  BUFX12 U1188 ( .A(n1807), .Y(n1812) );
  OR2X1 U1189 ( .A(n2322), .B(n2321), .Y(n2448) );
  BUFX20 U1191 ( .A(n1808), .Y(n1813) );
  BUFX12 U1195 ( .A(n1809), .Y(n1808) );
  OAI2BB1X1 U1723 ( .A0N(n3251), .A1N(n3116), .B0(n2588), .Y(n790) );
  MXI2X1 U1758 ( .A(n2446), .B(n3236), .S0(n3126), .Y(n801) );
  NOR2X1 U1759 ( .A(n2437), .B(n3127), .Y(n2335) );
  NOR2X1 U1761 ( .A(n1800), .B(n3127), .Y(n2333) );
  OAI2BB1X1 U1762 ( .A0N(n3130), .A1N(n3129), .B0(n3128), .Y(n818) );
  CLKINVX1 U1763 ( .A(n818), .Y(n636) );
  NAND3X1 U1764 ( .A(n2317), .B(n818), .C(n2484), .Y(n2318) );
  NAND2X1 U1765 ( .A(n3132), .B(n3131), .Y(n2459) );
  NOR3X1 U1766 ( .A(n3134), .B(n3122), .C(n3133), .Y(n2462) );
  NOR2X1 U1771 ( .A(n3136), .B(n3135), .Y(n2626) );
  NAND2X1 U1772 ( .A(n3138), .B(n3137), .Y(n1463) );
  NOR2X1 U1774 ( .A(n3119), .B(n3140), .Y(n1459) );
  OAI21XL U1777 ( .A0(n3142), .A1(n3141), .B0(n3122), .Y(n2463) );
  CLKINVX1 U1781 ( .A(n2632), .Y(n2617) );
  NOR2X1 U1782 ( .A(n3144), .B(n3143), .Y(n2632) );
  MXI2X1 U1783 ( .A(n3147), .B(n3146), .S0(n3145), .Y(n2609) );
  OAI22XL U1785 ( .A0(n3121), .A1(n3149), .B0(n3120), .B1(n3148), .Y(n1490) );
  AOI21X1 U1787 ( .A0(n1490), .A1(n2469), .B0(n3171), .Y(n1487) );
  NAND2X1 U1789 ( .A(n3120), .B(n3150), .Y(n2469) );
  MXI2X1 U1797 ( .A(n3203), .B(n3202), .S0(n1800), .Y(n2446) );
  MXI2X1 U1799 ( .A(n3197), .B(n3196), .S0(n1800), .Y(n2443) );
  CLKINVX1 U1802 ( .A(n799), .Y(n618) );
  INVX4 U1803 ( .A(n806), .Y(n625) );
  CLKINVX1 U1807 ( .A(n794), .Y(n613) );
  MXI2X1 U1808 ( .A(n2888), .B(n3183), .S0(n1800), .Y(n2442) );
  MXI2X1 U1810 ( .A(n2886), .B(n3175), .S0(n1800), .Y(n2436) );
  OAI2BB1X2 U1838 ( .A0N(n2881), .A1N(n2335), .B0(n2324), .Y(n802) );
  CLKINVX1 U1839 ( .A(n796), .Y(n615) );
  INVX3 U2076 ( .A(n3151), .Y(n1800) );
  MXI2X1 U2232 ( .A(n2885), .B(n3182), .S0(n1800), .Y(n2449) );
  MXI2X1 U2290 ( .A(n2887), .B(n3176), .S0(n1800), .Y(n2383) );
  NAND2X1 U2291 ( .A(n2626), .B(n3152), .Y(n1456) );
  OR2X1 U2293 ( .A(n3154), .B(n3153), .Y(n1454) );
  NOR2X1 U2294 ( .A(n2632), .B(n1463), .Y(n2635) );
  AND2X2 U2295 ( .A(n3156), .B(n3155), .Y(n993) );
  OR2X1 U2296 ( .A(n2632), .B(n3157), .Y(n1465) );
  OAI21XL U2297 ( .A0(n3160), .A1(n3159), .B0(n3158), .Y(n1447) );
  AOI22X1 U2298 ( .A0(n3164), .A1(n3163), .B0(n3162), .B1(n3161), .Y(n2380) );
  NAND3X1 U2299 ( .A(n2617), .B(n2618), .C(n1459), .Y(n1458) );
  AOI21X1 U2300 ( .A0(n3167), .A1(n3166), .B0(n3165), .Y(n2627) );
  NAND2X1 U2301 ( .A(n3169), .B(n3168), .Y(n2453) );
  OA21XL U2304 ( .A0(n2609), .A1(n3116), .B0(n1454), .Y(n996) );
  OR2X1 U2305 ( .A(n2626), .B(n3172), .Y(n2634) );
  MXI2X1 U2306 ( .A(n2437), .B(n3174), .S0(n3173), .Y(n810) );
  INVX3 U2308 ( .A(n1800), .Y(n2437) );
  CLKINVX1 U2329 ( .A(n810), .Y(n1726) );
  OA21XL U2337 ( .A0(n2609), .A1(n3117), .B0(n1454), .Y(n1136) );
  NAND3BX1 U2346 ( .AN(n3178), .B(n2459), .C(n3177), .Y(n2460) );
  OAI22XL U2347 ( .A0(n3123), .A1(n3181), .B0(n3180), .B1(n3179), .Y(n2470) );
  CLKINVX1 U2348 ( .A(n2635), .Y(n1462) );
  NAND3X1 U2349 ( .A(n2617), .B(n2618), .C(n3184), .Y(n1051) );
  MXI2X1 U2353 ( .A(n3186), .B(n3185), .S0(n2437), .Y(n2328) );
  OAI2BB1X1 U2457 ( .A0N(n3188), .A1N(n3187), .B0(n1447), .Y(n2475) );
  NAND2BX1 U2467 ( .AN(n2466), .B(n3189), .Y(n1491) );
  NAND2X1 U2471 ( .A(n2609), .B(n3117), .Y(n2610) );
  AOI21X1 U2473 ( .A0(n2463), .A1(n3192), .B0(n2462), .Y(n1101) );
  MXI2X1 U2474 ( .A(n3193), .B(n2877), .S0(n1800), .Y(n2325) );
  MXI2X1 U2481 ( .A(n3195), .B(n3194), .S0(n1800), .Y(n2444) );
  NOR2X1 U2483 ( .A(n1051), .B(n3198), .Y(n1050) );
  OAI22XL U2485 ( .A0(n2380), .A1(n3201), .B0(n3200), .B1(n3199), .Y(n2381) );
  AOI2BB2X1 U2501 ( .B0(n3205), .B1(n2333), .A0N(n3118), .A1N(n3204), .Y(n2334) );
  NAND3X1 U2502 ( .A(n2889), .B(n3206), .C(n2437), .Y(n2441) );
  OAI21XL U2503 ( .A0(n3207), .A1(n3115), .B0(n2460), .Y(n2464) );
  OAI31XL U2504 ( .A0(n1465), .A1(n3119), .A2(n3208), .B0(n1462), .Y(n1461) );
  NAND2X1 U2505 ( .A(n1458), .B(n1456), .Y(n1455) );
  OAI21XL U2506 ( .A0(n3210), .A1(n3209), .B0(n993), .Y(n1452) );
  NAND2X1 U2507 ( .A(N1215), .B(n3124), .Y(n2587) );
  MXI2X1 U2508 ( .A(n3212), .B(n3211), .S0(n2437), .Y(n2327) );
  CLKINVX1 U2509 ( .A(n2470), .Y(n1484) );
  OAI2BB1X1 U2510 ( .A0N(n3214), .A1N(n3213), .B0(n2458), .Y(n2465) );
  MXI2X1 U2511 ( .A(n3216), .B(n3215), .S0(n2437), .Y(n2329) );
  AOI2BB2X1 U2523 ( .B0(n3218), .B1(n2333), .A0N(n3118), .A1N(n3217), .Y(n2324) );
  NAND2X1 U2527 ( .A(n1491), .B(n3219), .Y(n1485) );
  NAND2X1 U2528 ( .A(n2475), .B(n3220), .Y(n2490) );
  NOR2BX1 U2541 ( .AN(n2627), .B(n1455), .Y(n2628) );
  NAND2X1 U2543 ( .A(N1216), .B(n3124), .Y(n1057) );
  OAI2BB1X1 U2545 ( .A0N(n3121), .A1N(n3221), .B0(n2453), .Y(n2456) );
  MXI2X1 U2547 ( .A(n2878), .B(n3222), .S0(n2437), .Y(n2326) );
  MXI2X1 U2549 ( .A(n2879), .B(n3223), .S0(n2437), .Y(n2331) );
  OAI21X1 U2559 ( .A0(n3125), .A1(n3224), .B0(n2587), .Y(n793) );
  CLKINVX1 U2580 ( .A(n793), .Y(n612) );
  MXI2X2 U2581 ( .A(n2436), .B(n3225), .S0(n3126), .Y(n797) );
  CLKINVX1 U2582 ( .A(n797), .Y(n616) );
  OAI2BB1X1 U2584 ( .A0N(n2335), .A1N(n2880), .B0(n2334), .Y(n803) );
  CLKINVX1 U2585 ( .A(n803), .Y(n622) );
  NOR3X1 U2589 ( .A(n2456), .B(n2455), .C(n2470), .Y(n2472) );
  OAI2BB1X1 U2684 ( .A0N(n1136), .A1N(n1452), .B0(n2610), .Y(n1066) );
  CLKINVX1 U2688 ( .A(n1050), .Y(n1049) );
  NAND2X1 U2689 ( .A(n1485), .B(n1484), .Y(n1483) );
  OAI2BB1X1 U2718 ( .A0N(n3226), .A1N(n2635), .B0(n2628), .Y(n2639) );
  CLKINVX1 U2722 ( .A(n802), .Y(n621) );
  NAND2X1 U2723 ( .A(N1217), .B(n3124), .Y(n2586) );
  OAI2BB1X1 U2724 ( .A0N(n2475), .A1N(n3228), .B0(n3227), .Y(n2382) );
  AND2X2 U2727 ( .A(n1491), .B(n1487), .Y(n1091) );
  NAND2X1 U2824 ( .A(n1057), .B(n3229), .Y(n792) );
  CLKINVX1 U2914 ( .A(n792), .Y(n611) );
  NAND2X1 U3250 ( .A(N1218), .B(n3124), .Y(n2588) );
  CLKINVX1 U3251 ( .A(n776), .Y(n1735) );
  AOI211XL U3252 ( .A0(n776), .A1(n2905), .B0(n2818), .C0(n2817), .Y(n2821) );
  MXI2X2 U3253 ( .A(n2444), .B(n3115), .S0(n3126), .Y(n799) );
  NAND3X1 U3254 ( .A(n2441), .B(n2440), .C(n3235), .Y(n794) );
  OAI21XL U3255 ( .A0(n2464), .A1(n2465), .B0(n1101), .Y(n2471) );
  CLKINVX1 U3256 ( .A(n801), .Y(n620) );
  AOI2BB2X1 U3332 ( .B0(n2381), .B1(n3239), .A0N(n3238), .A1N(n3237), .Y(n1144) );
  OAI2BB1X1 U3333 ( .A0N(n3125), .A1N(N1220), .B0(n3252), .Y(n2864) );
  NOR2X1 U3334 ( .A(n1461), .B(n2634), .Y(n2636) );
  OAI2BB1X1 U3335 ( .A0N(n996), .A1N(n1452), .B0(n2610), .Y(n2637) );
  CLKINVX1 U3336 ( .A(n800), .Y(n619) );
  CLKINVX1 U3337 ( .A(n795), .Y(n614) );
  INVX4 U3338 ( .A(n798), .Y(n617) );
  MXI2X2 U3339 ( .A(n2327), .B(n3243), .S0(n3127), .Y(n809) );
  CLKINVX1 U3340 ( .A(n809), .Y(n628) );
  INVX4 U3341 ( .A(n807), .Y(n626) );
  CLKINVX1 U3342 ( .A(n808), .Y(n627) );
  NOR2X1 U3343 ( .A(n2637), .B(n1049), .Y(n2640) );
  MXI2X2 U3344 ( .A(n2331), .B(n3247), .S0(n3127), .Y(n804) );
  CLKINVX1 U3345 ( .A(n804), .Y(n623) );
  OAI21X1 U3346 ( .A0(n3125), .A1(n3248), .B0(n2586), .Y(n791) );
  INVX3 U3347 ( .A(n791), .Y(n610) );
  NAND2X1 U3348 ( .A(n2382), .B(n1144), .Y(n782) );
  INVX3 U3349 ( .A(n782), .Y(n1116) );
  INVX4 U3350 ( .A(n805), .Y(n624) );
  OAI21XL U3351 ( .A0(n1066), .A1(n1051), .B0(n2636), .Y(n2638) );
  AOI2BB2X2 U3352 ( .B0(n2472), .B1(n2471), .A0N(n1091), .A1N(n1483), .Y(n775)
         );
  CLKINVX1 U3353 ( .A(n775), .Y(n1719) );
  OAI2BB1X1 U3354 ( .A0N(n3125), .A1N(N1219), .B0(n3250), .Y(n2861) );
  CLKINVX1 U3355 ( .A(n2861), .Y(n608) );
  NAND2X4 U3356 ( .A(n2630), .B(n2861), .Y(n2616) );
  OAI21X1 U3357 ( .A0(n2640), .A1(n2639), .B0(n2638), .Y(n2865) );
  CLKINVX1 U3358 ( .A(n2865), .Y(n1742) );
  INVX4 U3359 ( .A(n2864), .Y(n607) );
  OAI2BB1X1 U3360 ( .A0N(n3125), .A1N(N1222), .B0(n3253), .Y(n2862) );
  CLKINVX1 U3361 ( .A(n2862), .Y(n605) );
  OAI2BB1X1 U3362 ( .A0N(n3125), .A1N(N1221), .B0(n3254), .Y(n2863) );
  CLKINVX1 U3363 ( .A(n2863), .Y(n606) );
endmodule

